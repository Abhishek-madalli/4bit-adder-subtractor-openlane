magic
tech sky130A
magscale 1 2
timestamp 1755103505
<< viali >>
rect 1593 10761 1627 10795
rect 1501 10625 1535 10659
rect 1961 10625 1995 10659
rect 4169 10625 4203 10659
rect 4629 10625 4663 10659
rect 4813 10625 4847 10659
rect 4905 10625 4939 10659
rect 5273 10625 5307 10659
rect 5457 10625 5491 10659
rect 7389 10625 7423 10659
rect 9505 10625 9539 10659
rect 9781 10625 9815 10659
rect 2145 10421 2179 10455
rect 3985 10421 4019 10455
rect 4445 10421 4479 10455
rect 5089 10421 5123 10455
rect 7205 10421 7239 10455
rect 9321 10421 9355 10455
rect 9597 10421 9631 10455
rect 2126 10217 2160 10251
rect 3617 10217 3651 10251
rect 5089 10217 5123 10251
rect 6579 10217 6613 10251
rect 1869 10081 1903 10115
rect 4445 10081 4479 10115
rect 6837 10081 6871 10115
rect 6929 10081 6963 10115
rect 7205 10081 7239 10115
rect 4537 10013 4571 10047
rect 4813 10013 4847 10047
rect 4997 10013 5031 10047
rect 4169 9877 4203 9911
rect 4997 9877 5031 9911
rect 8677 9877 8711 9911
rect 1409 9673 1443 9707
rect 4445 9673 4479 9707
rect 4905 9673 4939 9707
rect 5625 9673 5659 9707
rect 2881 9605 2915 9639
rect 5825 9605 5859 9639
rect 4353 9537 4387 9571
rect 4629 9537 4663 9571
rect 5365 9537 5399 9571
rect 3157 9469 3191 9503
rect 4813 9333 4847 9367
rect 5273 9333 5307 9367
rect 5457 9333 5491 9367
rect 5641 9333 5675 9367
rect 7021 8925 7055 8959
rect 9781 8925 9815 8959
rect 1501 8857 1535 8891
rect 1593 8789 1627 8823
rect 6469 8789 6503 8823
rect 9597 8789 9631 8823
rect 1409 8585 1443 8619
rect 3709 8517 3743 8551
rect 5549 8517 5583 8551
rect 8125 8517 8159 8551
rect 5365 8449 5399 8483
rect 2881 8381 2915 8415
rect 3157 8381 3191 8415
rect 3433 8381 3467 8415
rect 8401 8381 8435 8415
rect 6653 8313 6687 8347
rect 5181 8245 5215 8279
rect 5457 7905 5491 7939
rect 5733 7905 5767 7939
rect 6009 7905 6043 7939
rect 6561 7905 6595 7939
rect 5365 7837 5399 7871
rect 6101 7837 6135 7871
rect 5273 7769 5307 7803
rect 6837 7769 6871 7803
rect 4905 7701 4939 7735
rect 8309 7701 8343 7735
rect 3065 7497 3099 7531
rect 4445 7497 4479 7531
rect 5549 7497 5583 7531
rect 4353 7361 4387 7395
rect 4813 7361 4847 7395
rect 5089 7361 5123 7395
rect 5181 7361 5215 7395
rect 5365 7361 5399 7395
rect 8401 7361 8435 7395
rect 4905 7293 4939 7327
rect 9045 7157 9079 7191
rect 4997 6953 5031 6987
rect 4629 6817 4663 6851
rect 6745 6817 6779 6851
rect 5089 6749 5123 6783
rect 5181 6681 5215 6715
rect 4629 6409 4663 6443
rect 5549 6409 5583 6443
rect 8486 6409 8520 6443
rect 4353 6341 4387 6375
rect 4537 6341 4571 6375
rect 4997 6341 5031 6375
rect 5181 6341 5215 6375
rect 5381 6341 5415 6375
rect 8017 6341 8051 6375
rect 8217 6341 8251 6375
rect 8585 6341 8619 6375
rect 4169 6273 4203 6307
rect 4813 6273 4847 6307
rect 5089 6273 5123 6307
rect 7481 6273 7515 6307
rect 7665 6273 7699 6307
rect 8309 6273 8343 6307
rect 8401 6273 8435 6307
rect 7849 6137 7883 6171
rect 5365 6069 5399 6103
rect 7665 6069 7699 6103
rect 8033 6069 8067 6103
rect 4813 5865 4847 5899
rect 9045 5865 9079 5899
rect 5641 5729 5675 5763
rect 1409 5661 1443 5695
rect 4169 5661 4203 5695
rect 4721 5661 4755 5695
rect 4905 5661 4939 5695
rect 7021 5661 7055 5695
rect 8953 5661 8987 5695
rect 9137 5661 9171 5695
rect 7297 5593 7331 5627
rect 9413 5593 9447 5627
rect 1593 5525 1627 5559
rect 4077 5525 4111 5559
rect 4997 5525 5031 5559
rect 8769 5525 8803 5559
rect 9689 5525 9723 5559
rect 1869 5321 1903 5355
rect 7021 5321 7055 5355
rect 8217 5321 8251 5355
rect 5181 5253 5215 5287
rect 8401 5253 8435 5287
rect 6653 5185 6687 5219
rect 7205 5185 7239 5219
rect 7297 5185 7331 5219
rect 7573 5185 7607 5219
rect 7849 5185 7883 5219
rect 8033 5185 8067 5219
rect 8585 5185 8619 5219
rect 3341 5117 3375 5151
rect 3617 5117 3651 5151
rect 3709 5117 3743 5151
rect 5457 5117 5491 5151
rect 6929 5117 6963 5151
rect 7481 5117 7515 5151
rect 8125 5117 8159 5151
rect 6469 4981 6503 5015
rect 6837 4981 6871 5015
rect 7665 4981 7699 5015
rect 7205 4777 7239 4811
rect 7573 4777 7607 4811
rect 7113 4573 7147 4607
rect 7297 4573 7331 4607
rect 7665 4573 7699 4607
rect 7297 3553 7331 3587
rect 7021 3485 7055 3519
rect 8769 3349 8803 3383
rect 8585 3145 8619 3179
rect 3709 3077 3743 3111
rect 5273 3077 5307 3111
rect 1501 3009 1535 3043
rect 9505 3009 9539 3043
rect 3801 2941 3835 2975
rect 5549 2941 5583 2975
rect 6837 2941 6871 2975
rect 7113 2941 7147 2975
rect 1593 2805 1627 2839
rect 2421 2805 2455 2839
rect 9689 2805 9723 2839
rect 1409 2601 1443 2635
rect 3249 2601 3283 2635
rect 8493 2601 8527 2635
rect 9597 2601 9631 2635
rect 3157 2465 3191 2499
rect 3433 2397 3467 2431
rect 5181 2397 5215 2431
rect 8677 2397 8711 2431
rect 9781 2397 9815 2431
rect 2881 2329 2915 2363
rect 5273 2261 5307 2295
<< metal1 >>
rect 1104 10906 10120 10928
rect 1104 10854 2737 10906
rect 2789 10854 2801 10906
rect 2853 10854 2865 10906
rect 2917 10854 2929 10906
rect 2981 10854 2993 10906
rect 3045 10854 4991 10906
rect 5043 10854 5055 10906
rect 5107 10854 5119 10906
rect 5171 10854 5183 10906
rect 5235 10854 5247 10906
rect 5299 10854 7245 10906
rect 7297 10854 7309 10906
rect 7361 10854 7373 10906
rect 7425 10854 7437 10906
rect 7489 10854 7501 10906
rect 7553 10854 9499 10906
rect 9551 10854 9563 10906
rect 9615 10854 9627 10906
rect 9679 10854 9691 10906
rect 9743 10854 9755 10906
rect 9807 10854 10120 10906
rect 1104 10832 10120 10854
rect 1302 10752 1308 10804
rect 1360 10792 1366 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1360 10764 1593 10792
rect 1360 10752 1366 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 7098 10752 7104 10804
rect 7156 10752 7162 10804
rect 9306 10752 9312 10804
rect 9364 10752 9370 10804
rect 9858 10752 9864 10804
rect 9916 10752 9922 10804
rect 4632 10696 5856 10724
rect 1486 10616 1492 10668
rect 1544 10616 1550 10668
rect 1946 10616 1952 10668
rect 2004 10616 2010 10668
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 4632 10665 4660 10696
rect 5828 10668 5856 10696
rect 4157 10659 4215 10665
rect 4157 10656 4169 10659
rect 3936 10628 4169 10656
rect 3936 10616 3942 10628
rect 4157 10625 4169 10628
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 4801 10659 4859 10665
rect 4801 10625 4813 10659
rect 4847 10625 4859 10659
rect 4801 10619 4859 10625
rect 4893 10659 4951 10665
rect 4893 10625 4905 10659
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 3602 10548 3608 10600
rect 3660 10588 3666 10600
rect 4632 10588 4660 10619
rect 3660 10560 4660 10588
rect 3660 10548 3666 10560
rect 4816 10520 4844 10619
rect 4908 10588 4936 10619
rect 5258 10616 5264 10668
rect 5316 10616 5322 10668
rect 5442 10616 5448 10668
rect 5500 10616 5506 10668
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 7116 10656 7144 10752
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 7116 10628 7389 10656
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 9324 10656 9352 10752
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 9324 10628 9505 10656
rect 7377 10619 7435 10625
rect 9493 10625 9505 10628
rect 9539 10625 9551 10659
rect 9493 10619 9551 10625
rect 9769 10659 9827 10665
rect 9769 10625 9781 10659
rect 9815 10656 9827 10659
rect 9876 10656 9904 10752
rect 9815 10628 9904 10656
rect 9815 10625 9827 10628
rect 9769 10619 9827 10625
rect 4908 10560 5672 10588
rect 4816 10492 5120 10520
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 2133 10455 2191 10461
rect 2133 10452 2145 10455
rect 2004 10424 2145 10452
rect 2004 10412 2010 10424
rect 2133 10421 2145 10424
rect 2179 10421 2191 10455
rect 2133 10415 2191 10421
rect 3970 10412 3976 10464
rect 4028 10412 4034 10464
rect 4246 10412 4252 10464
rect 4304 10452 4310 10464
rect 5092 10461 5120 10492
rect 5644 10464 5672 10560
rect 4433 10455 4491 10461
rect 4433 10452 4445 10455
rect 4304 10424 4445 10452
rect 4304 10412 4310 10424
rect 4433 10421 4445 10424
rect 4479 10421 4491 10455
rect 4433 10415 4491 10421
rect 5077 10455 5135 10461
rect 5077 10421 5089 10455
rect 5123 10452 5135 10455
rect 5534 10452 5540 10464
rect 5123 10424 5540 10452
rect 5123 10421 5135 10424
rect 5077 10415 5135 10421
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 5626 10412 5632 10464
rect 5684 10412 5690 10464
rect 6362 10412 6368 10464
rect 6420 10452 6426 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 6420 10424 7205 10452
rect 6420 10412 6426 10424
rect 7193 10421 7205 10424
rect 7239 10421 7251 10455
rect 7193 10415 7251 10421
rect 9306 10412 9312 10464
rect 9364 10412 9370 10464
rect 9582 10412 9588 10464
rect 9640 10412 9646 10464
rect 1104 10362 10120 10384
rect 1104 10310 2077 10362
rect 2129 10310 2141 10362
rect 2193 10310 2205 10362
rect 2257 10310 2269 10362
rect 2321 10310 2333 10362
rect 2385 10310 4331 10362
rect 4383 10310 4395 10362
rect 4447 10310 4459 10362
rect 4511 10310 4523 10362
rect 4575 10310 4587 10362
rect 4639 10310 6585 10362
rect 6637 10310 6649 10362
rect 6701 10310 6713 10362
rect 6765 10310 6777 10362
rect 6829 10310 6841 10362
rect 6893 10310 8839 10362
rect 8891 10310 8903 10362
rect 8955 10310 8967 10362
rect 9019 10310 9031 10362
rect 9083 10310 9095 10362
rect 9147 10310 10120 10362
rect 1104 10288 10120 10310
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 2114 10251 2172 10257
rect 2114 10248 2126 10251
rect 2004 10220 2126 10248
rect 2004 10208 2010 10220
rect 2114 10217 2126 10220
rect 2160 10217 2172 10251
rect 2114 10211 2172 10217
rect 3602 10208 3608 10260
rect 3660 10208 3666 10260
rect 5077 10251 5135 10257
rect 5077 10217 5089 10251
rect 5123 10248 5135 10251
rect 5258 10248 5264 10260
rect 5123 10220 5264 10248
rect 5123 10217 5135 10220
rect 5077 10211 5135 10217
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 6567 10251 6625 10257
rect 6567 10217 6579 10251
rect 6613 10248 6625 10251
rect 9306 10248 9312 10260
rect 6613 10220 9312 10248
rect 6613 10217 6625 10220
rect 6567 10211 6625 10217
rect 9306 10208 9312 10220
rect 9364 10208 9370 10260
rect 9582 10208 9588 10260
rect 9640 10208 9646 10260
rect 1857 10115 1915 10121
rect 1857 10081 1869 10115
rect 1903 10112 1915 10115
rect 3418 10112 3424 10124
rect 1903 10084 3424 10112
rect 1903 10081 1915 10084
rect 1857 10075 1915 10081
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 4430 10072 4436 10124
rect 4488 10072 4494 10124
rect 5166 10112 5172 10124
rect 4816 10084 5172 10112
rect 4522 10004 4528 10056
rect 4580 10004 4586 10056
rect 4816 10053 4844 10084
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 5258 10072 5264 10124
rect 5316 10072 5322 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6825 10115 6883 10121
rect 6825 10112 6837 10115
rect 6512 10084 6837 10112
rect 6512 10072 6518 10084
rect 6825 10081 6837 10084
rect 6871 10112 6883 10115
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 6871 10084 6929 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 6917 10081 6929 10084
rect 6963 10081 6975 10115
rect 6917 10075 6975 10081
rect 7193 10115 7251 10121
rect 7193 10081 7205 10115
rect 7239 10112 7251 10115
rect 9600 10112 9628 10208
rect 7239 10084 9628 10112
rect 7239 10081 7251 10084
rect 7193 10075 7251 10081
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10044 5043 10047
rect 5276 10044 5304 10072
rect 5031 10016 5304 10044
rect 5031 10013 5043 10016
rect 4985 10007 5043 10013
rect 4706 9976 4712 9988
rect 3358 9948 4712 9976
rect 4706 9936 4712 9948
rect 4764 9976 4770 9988
rect 4764 9948 5382 9976
rect 4764 9936 4770 9948
rect 7098 9936 7104 9988
rect 7156 9976 7162 9988
rect 7156 9948 7682 9976
rect 7156 9936 7162 9948
rect 4154 9868 4160 9920
rect 4212 9868 4218 9920
rect 4985 9911 5043 9917
rect 4985 9877 4997 9911
rect 5031 9908 5043 9911
rect 5626 9908 5632 9920
rect 5031 9880 5632 9908
rect 5031 9877 5043 9880
rect 4985 9871 5043 9877
rect 5626 9868 5632 9880
rect 5684 9868 5690 9920
rect 8662 9868 8668 9920
rect 8720 9868 8726 9920
rect 1104 9818 10120 9840
rect 1104 9766 2737 9818
rect 2789 9766 2801 9818
rect 2853 9766 2865 9818
rect 2917 9766 2929 9818
rect 2981 9766 2993 9818
rect 3045 9766 4991 9818
rect 5043 9766 5055 9818
rect 5107 9766 5119 9818
rect 5171 9766 5183 9818
rect 5235 9766 5247 9818
rect 5299 9766 7245 9818
rect 7297 9766 7309 9818
rect 7361 9766 7373 9818
rect 7425 9766 7437 9818
rect 7489 9766 7501 9818
rect 7553 9766 9499 9818
rect 9551 9766 9563 9818
rect 9615 9766 9627 9818
rect 9679 9766 9691 9818
rect 9743 9766 9755 9818
rect 9807 9766 10120 9818
rect 1104 9744 10120 9766
rect 1397 9707 1455 9713
rect 1397 9673 1409 9707
rect 1443 9704 1455 9707
rect 1486 9704 1492 9716
rect 1443 9676 1492 9704
rect 1443 9673 1455 9676
rect 1397 9667 1455 9673
rect 1486 9664 1492 9676
rect 1544 9664 1550 9716
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4433 9707 4491 9713
rect 4433 9704 4445 9707
rect 4304 9676 4445 9704
rect 4304 9664 4310 9676
rect 4433 9673 4445 9676
rect 4479 9673 4491 9707
rect 4433 9667 4491 9673
rect 2869 9639 2927 9645
rect 2869 9605 2881 9639
rect 2915 9636 2927 9639
rect 4154 9636 4160 9648
rect 2915 9608 4160 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 4448 9636 4476 9667
rect 4522 9664 4528 9716
rect 4580 9704 4586 9716
rect 5626 9713 5632 9716
rect 4893 9707 4951 9713
rect 4893 9704 4905 9707
rect 4580 9676 4905 9704
rect 4580 9664 4586 9676
rect 4893 9673 4905 9676
rect 4939 9673 4951 9707
rect 4893 9667 4951 9673
rect 5613 9707 5632 9713
rect 5613 9673 5625 9707
rect 5613 9667 5632 9673
rect 5626 9664 5632 9667
rect 5684 9664 5690 9716
rect 4448 9608 5396 9636
rect 5368 9577 5396 9608
rect 5810 9596 5816 9648
rect 5868 9596 5874 9648
rect 4341 9571 4399 9577
rect 1780 9500 1808 9554
rect 4341 9537 4353 9571
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 5353 9571 5411 9577
rect 4663 9540 5304 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 3145 9503 3203 9509
rect 1780 9472 3096 9500
rect 3068 9364 3096 9472
rect 3145 9469 3157 9503
rect 3191 9500 3203 9503
rect 3418 9500 3424 9512
rect 3191 9472 3424 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 4356 9500 4384 9531
rect 4430 9500 4436 9512
rect 4356 9472 4436 9500
rect 4430 9460 4436 9472
rect 4488 9500 4494 9512
rect 4488 9472 5212 9500
rect 4488 9460 4494 9472
rect 5184 9376 5212 9472
rect 3234 9364 3240 9376
rect 3068 9336 3240 9364
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 4798 9324 4804 9376
rect 4856 9324 4862 9376
rect 5166 9324 5172 9376
rect 5224 9324 5230 9376
rect 5276 9373 5304 9540
rect 5353 9537 5365 9571
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5261 9367 5319 9373
rect 5261 9333 5273 9367
rect 5307 9364 5319 9367
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 5307 9336 5457 9364
rect 5307 9333 5319 9336
rect 5261 9327 5319 9333
rect 5445 9333 5457 9336
rect 5491 9333 5503 9367
rect 5445 9327 5503 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 5629 9367 5687 9373
rect 5629 9364 5641 9367
rect 5592 9336 5641 9364
rect 5592 9324 5598 9336
rect 5629 9333 5641 9336
rect 5675 9333 5687 9367
rect 5629 9327 5687 9333
rect 1104 9274 10120 9296
rect 1104 9222 2077 9274
rect 2129 9222 2141 9274
rect 2193 9222 2205 9274
rect 2257 9222 2269 9274
rect 2321 9222 2333 9274
rect 2385 9222 4331 9274
rect 4383 9222 4395 9274
rect 4447 9222 4459 9274
rect 4511 9222 4523 9274
rect 4575 9222 4587 9274
rect 4639 9222 6585 9274
rect 6637 9222 6649 9274
rect 6701 9222 6713 9274
rect 6765 9222 6777 9274
rect 6829 9222 6841 9274
rect 6893 9222 8839 9274
rect 8891 9222 8903 9274
rect 8955 9222 8967 9274
rect 9019 9222 9031 9274
rect 9083 9222 9095 9274
rect 9147 9222 10120 9274
rect 1104 9200 10120 9222
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 6914 9160 6920 9172
rect 4856 9132 6920 9160
rect 4856 9120 4862 9132
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 7009 8959 7067 8965
rect 7009 8956 7021 8959
rect 6696 8928 7021 8956
rect 6696 8916 6702 8928
rect 7009 8925 7021 8928
rect 7055 8925 7067 8959
rect 7009 8919 7067 8925
rect 9769 8959 9827 8965
rect 9769 8925 9781 8959
rect 9815 8956 9827 8959
rect 10134 8956 10140 8968
rect 9815 8928 10140 8956
rect 9815 8925 9827 8928
rect 9769 8919 9827 8925
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 1486 8848 1492 8900
rect 1544 8848 1550 8900
rect 934 8780 940 8832
rect 992 8820 998 8832
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 992 8792 1593 8820
rect 992 8780 998 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 6270 8780 6276 8832
rect 6328 8820 6334 8832
rect 6457 8823 6515 8829
rect 6457 8820 6469 8823
rect 6328 8792 6469 8820
rect 6328 8780 6334 8792
rect 6457 8789 6469 8792
rect 6503 8789 6515 8823
rect 6457 8783 6515 8789
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9585 8823 9643 8829
rect 9585 8820 9597 8823
rect 8904 8792 9597 8820
rect 8904 8780 8910 8792
rect 9585 8789 9597 8792
rect 9631 8789 9643 8823
rect 9585 8783 9643 8789
rect 1104 8730 10120 8752
rect 1104 8678 2737 8730
rect 2789 8678 2801 8730
rect 2853 8678 2865 8730
rect 2917 8678 2929 8730
rect 2981 8678 2993 8730
rect 3045 8678 4991 8730
rect 5043 8678 5055 8730
rect 5107 8678 5119 8730
rect 5171 8678 5183 8730
rect 5235 8678 5247 8730
rect 5299 8678 7245 8730
rect 7297 8678 7309 8730
rect 7361 8678 7373 8730
rect 7425 8678 7437 8730
rect 7489 8678 7501 8730
rect 7553 8678 9499 8730
rect 9551 8678 9563 8730
rect 9615 8678 9627 8730
rect 9679 8678 9691 8730
rect 9743 8678 9755 8730
rect 9807 8678 10120 8730
rect 1104 8656 10120 8678
rect 1397 8619 1455 8625
rect 1397 8585 1409 8619
rect 1443 8616 1455 8619
rect 1486 8616 1492 8628
rect 1443 8588 1492 8616
rect 1443 8585 1455 8588
rect 1397 8579 1455 8585
rect 1486 8576 1492 8588
rect 1544 8576 1550 8628
rect 4706 8576 4712 8628
rect 4764 8616 4770 8628
rect 7098 8616 7104 8628
rect 4764 8588 5028 8616
rect 4764 8576 4770 8588
rect 3234 8548 3240 8560
rect 2438 8520 3240 8548
rect 3234 8508 3240 8520
rect 3292 8508 3298 8560
rect 3697 8551 3755 8557
rect 3697 8517 3709 8551
rect 3743 8548 3755 8551
rect 3970 8548 3976 8560
rect 3743 8520 3976 8548
rect 3743 8517 3755 8520
rect 3697 8511 3755 8517
rect 3970 8508 3976 8520
rect 4028 8508 4034 8560
rect 5000 8548 5028 8588
rect 5552 8588 7104 8616
rect 5552 8557 5580 8588
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 8202 8616 8208 8628
rect 7760 8588 8208 8616
rect 5537 8551 5595 8557
rect 5537 8548 5549 8551
rect 4922 8520 5549 8548
rect 5537 8517 5549 8520
rect 5583 8517 5595 8551
rect 7760 8548 7788 8588
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 8846 8576 8852 8628
rect 8904 8576 8910 8628
rect 7682 8520 7788 8548
rect 8113 8551 8171 8557
rect 5537 8511 5595 8517
rect 8113 8517 8125 8551
rect 8159 8548 8171 8551
rect 8864 8548 8892 8576
rect 8159 8520 8892 8548
rect 8159 8517 8171 8520
rect 8113 8511 8171 8517
rect 5353 8483 5411 8489
rect 5353 8449 5365 8483
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8412 2927 8415
rect 3145 8415 3203 8421
rect 2915 8384 3096 8412
rect 2915 8381 2927 8384
rect 2869 8375 2927 8381
rect 3068 8344 3096 8384
rect 3145 8381 3157 8415
rect 3191 8412 3203 8415
rect 3418 8412 3424 8424
rect 3191 8384 3424 8412
rect 3191 8381 3203 8384
rect 3145 8375 3203 8381
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 4154 8412 4160 8424
rect 3528 8384 4160 8412
rect 3528 8344 3556 8384
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 4706 8372 4712 8424
rect 4764 8412 4770 8424
rect 5368 8412 5396 8443
rect 4764 8384 5396 8412
rect 4764 8372 4770 8384
rect 8386 8372 8392 8424
rect 8444 8372 8450 8424
rect 3068 8316 3556 8344
rect 6638 8304 6644 8356
rect 6696 8304 6702 8356
rect 5166 8236 5172 8288
rect 5224 8236 5230 8288
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 6656 8276 6684 8304
rect 5960 8248 6684 8276
rect 5960 8236 5966 8248
rect 1104 8186 10120 8208
rect 1104 8134 2077 8186
rect 2129 8134 2141 8186
rect 2193 8134 2205 8186
rect 2257 8134 2269 8186
rect 2321 8134 2333 8186
rect 2385 8134 4331 8186
rect 4383 8134 4395 8186
rect 4447 8134 4459 8186
rect 4511 8134 4523 8186
rect 4575 8134 4587 8186
rect 4639 8134 6585 8186
rect 6637 8134 6649 8186
rect 6701 8134 6713 8186
rect 6765 8134 6777 8186
rect 6829 8134 6841 8186
rect 6893 8134 8839 8186
rect 8891 8134 8903 8186
rect 8955 8134 8967 8186
rect 9019 8134 9031 8186
rect 9083 8134 9095 8186
rect 9147 8134 10120 8186
rect 1104 8112 10120 8134
rect 3418 8032 3424 8084
rect 3476 8072 3482 8084
rect 6454 8072 6460 8084
rect 3476 8044 6460 8072
rect 3476 8032 3482 8044
rect 6454 8032 6460 8044
rect 6512 8072 6518 8084
rect 8386 8072 8392 8084
rect 6512 8044 8392 8072
rect 6512 8032 6518 8044
rect 5460 7976 6040 8004
rect 5166 7896 5172 7948
rect 5224 7936 5230 7948
rect 5460 7945 5488 7976
rect 5445 7939 5503 7945
rect 5445 7936 5457 7939
rect 5224 7908 5457 7936
rect 5224 7896 5230 7908
rect 5445 7905 5457 7908
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 5718 7896 5724 7948
rect 5776 7896 5782 7948
rect 6012 7945 6040 7976
rect 6564 7945 6592 8044
rect 8386 8032 8392 8044
rect 8444 8032 8450 8084
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 6549 7939 6607 7945
rect 6549 7905 6561 7939
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7868 5411 7871
rect 5902 7868 5908 7880
rect 5399 7840 5908 7868
rect 5399 7837 5411 7840
rect 5353 7831 5411 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6270 7868 6276 7880
rect 6135 7840 6276 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 4246 7760 4252 7812
rect 4304 7800 4310 7812
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 4304 7772 5273 7800
rect 4304 7760 4310 7772
rect 5261 7769 5273 7772
rect 5307 7800 5319 7803
rect 5442 7800 5448 7812
rect 5307 7772 5448 7800
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 5442 7760 5448 7772
rect 5500 7760 5506 7812
rect 6362 7760 6368 7812
rect 6420 7800 6426 7812
rect 6825 7803 6883 7809
rect 6825 7800 6837 7803
rect 6420 7772 6837 7800
rect 6420 7760 6426 7772
rect 6825 7769 6837 7772
rect 6871 7769 6883 7803
rect 6825 7763 6883 7769
rect 7098 7760 7104 7812
rect 7156 7800 7162 7812
rect 7156 7772 7314 7800
rect 7156 7760 7162 7772
rect 4890 7692 4896 7744
rect 4948 7692 4954 7744
rect 8294 7692 8300 7744
rect 8352 7692 8358 7744
rect 1104 7642 10120 7664
rect 1104 7590 2737 7642
rect 2789 7590 2801 7642
rect 2853 7590 2865 7642
rect 2917 7590 2929 7642
rect 2981 7590 2993 7642
rect 3045 7590 4991 7642
rect 5043 7590 5055 7642
rect 5107 7590 5119 7642
rect 5171 7590 5183 7642
rect 5235 7590 5247 7642
rect 5299 7590 7245 7642
rect 7297 7590 7309 7642
rect 7361 7590 7373 7642
rect 7425 7590 7437 7642
rect 7489 7590 7501 7642
rect 7553 7590 9499 7642
rect 9551 7590 9563 7642
rect 9615 7590 9627 7642
rect 9679 7590 9691 7642
rect 9743 7590 9755 7642
rect 9807 7590 10120 7642
rect 1104 7568 10120 7590
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3418 7528 3424 7540
rect 3099 7500 3424 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3418 7488 3424 7500
rect 3476 7488 3482 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4433 7531 4491 7537
rect 4433 7528 4445 7531
rect 4212 7500 4445 7528
rect 4212 7488 4218 7500
rect 4433 7497 4445 7500
rect 4479 7497 4491 7531
rect 4433 7491 4491 7497
rect 4890 7488 4896 7540
rect 4948 7488 4954 7540
rect 5350 7488 5356 7540
rect 5408 7528 5414 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 5408 7500 5549 7528
rect 5408 7488 5414 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 5537 7491 5595 7497
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4341 7395 4399 7401
rect 4341 7392 4353 7395
rect 4212 7364 4353 7392
rect 4212 7352 4218 7364
rect 4341 7361 4353 7364
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4798 7352 4804 7404
rect 4856 7352 4862 7404
rect 4908 7392 4936 7488
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4908 7364 5089 7392
rect 4908 7333 4936 7364
rect 5077 7361 5089 7364
rect 5123 7361 5135 7395
rect 5077 7355 5135 7361
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 5534 7392 5540 7404
rect 5399 7364 5540 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7293 4951 7327
rect 4893 7287 4951 7293
rect 5184 7256 5212 7355
rect 5534 7352 5540 7364
rect 5592 7352 5598 7404
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 8352 7364 8401 7392
rect 8352 7352 8358 7364
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 4908 7228 5212 7256
rect 4908 7200 4936 7228
rect 4890 7148 4896 7200
rect 4948 7148 4954 7200
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 9033 7191 9091 7197
rect 9033 7188 9045 7191
rect 8812 7160 9045 7188
rect 8812 7148 8818 7160
rect 9033 7157 9045 7160
rect 9079 7157 9091 7191
rect 9033 7151 9091 7157
rect 1104 7098 10120 7120
rect 1104 7046 2077 7098
rect 2129 7046 2141 7098
rect 2193 7046 2205 7098
rect 2257 7046 2269 7098
rect 2321 7046 2333 7098
rect 2385 7046 4331 7098
rect 4383 7046 4395 7098
rect 4447 7046 4459 7098
rect 4511 7046 4523 7098
rect 4575 7046 4587 7098
rect 4639 7046 6585 7098
rect 6637 7046 6649 7098
rect 6701 7046 6713 7098
rect 6765 7046 6777 7098
rect 6829 7046 6841 7098
rect 6893 7046 8839 7098
rect 8891 7046 8903 7098
rect 8955 7046 8967 7098
rect 9019 7046 9031 7098
rect 9083 7046 9095 7098
rect 9147 7046 10120 7098
rect 1104 7024 10120 7046
rect 4154 6944 4160 6996
rect 4212 6944 4218 6996
rect 4985 6987 5043 6993
rect 4985 6953 4997 6987
rect 5031 6984 5043 6987
rect 5534 6984 5540 6996
rect 5031 6956 5540 6984
rect 5031 6953 5043 6956
rect 4985 6947 5043 6953
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 4172 6916 4200 6944
rect 4172 6888 5580 6916
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 4798 6848 4804 6860
rect 4663 6820 4804 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 5552 6848 5580 6888
rect 6733 6851 6791 6857
rect 6733 6848 6745 6851
rect 5552 6820 6745 6848
rect 6733 6817 6745 6820
rect 6779 6817 6791 6851
rect 6733 6811 6791 6817
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4948 6752 5089 6780
rect 4948 6740 4954 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 5169 6715 5227 6721
rect 5169 6712 5181 6715
rect 4212 6684 5181 6712
rect 4212 6672 4218 6684
rect 5169 6681 5181 6684
rect 5215 6681 5227 6715
rect 5169 6675 5227 6681
rect 1104 6554 10120 6576
rect 1104 6502 2737 6554
rect 2789 6502 2801 6554
rect 2853 6502 2865 6554
rect 2917 6502 2929 6554
rect 2981 6502 2993 6554
rect 3045 6502 4991 6554
rect 5043 6502 5055 6554
rect 5107 6502 5119 6554
rect 5171 6502 5183 6554
rect 5235 6502 5247 6554
rect 5299 6502 7245 6554
rect 7297 6502 7309 6554
rect 7361 6502 7373 6554
rect 7425 6502 7437 6554
rect 7489 6502 7501 6554
rect 7553 6502 9499 6554
rect 9551 6502 9563 6554
rect 9615 6502 9627 6554
rect 9679 6502 9691 6554
rect 9743 6502 9755 6554
rect 9807 6502 10120 6554
rect 1104 6480 10120 6502
rect 4246 6400 4252 6452
rect 4304 6400 4310 6452
rect 4617 6443 4675 6449
rect 4617 6409 4629 6443
rect 4663 6440 4675 6443
rect 4890 6440 4896 6452
rect 4663 6412 4896 6440
rect 4663 6409 4675 6412
rect 4617 6403 4675 6409
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5074 6400 5080 6452
rect 5132 6400 5138 6452
rect 5534 6400 5540 6452
rect 5592 6400 5598 6452
rect 8474 6443 8532 6449
rect 8474 6440 8486 6443
rect 7852 6412 8486 6440
rect 4264 6372 4292 6400
rect 4341 6375 4399 6381
rect 4341 6372 4353 6375
rect 4264 6344 4353 6372
rect 4341 6341 4353 6344
rect 4387 6341 4399 6375
rect 4341 6335 4399 6341
rect 4525 6375 4583 6381
rect 4525 6341 4537 6375
rect 4571 6372 4583 6375
rect 4985 6375 5043 6381
rect 4985 6372 4997 6375
rect 4571 6344 4997 6372
rect 4571 6341 4583 6344
rect 4525 6335 4583 6341
rect 4985 6341 4997 6344
rect 5031 6341 5043 6375
rect 5092 6372 5120 6400
rect 5169 6375 5227 6381
rect 5169 6372 5181 6375
rect 5092 6344 5181 6372
rect 4985 6335 5043 6341
rect 5169 6341 5181 6344
rect 5215 6341 5227 6375
rect 5369 6375 5427 6381
rect 5369 6372 5381 6375
rect 5169 6335 5227 6341
rect 5276 6344 5381 6372
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4246 6304 4252 6316
rect 4203 6276 4252 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4356 6236 4384 6335
rect 4798 6264 4804 6316
rect 4856 6264 4862 6316
rect 4890 6236 4896 6248
rect 4356 6208 4896 6236
rect 4890 6196 4896 6208
rect 4948 6196 4954 6248
rect 5000 6100 5028 6335
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5276 6304 5304 6344
rect 5369 6341 5381 6344
rect 5415 6341 5427 6375
rect 5369 6335 5427 6341
rect 7852 6316 7880 6412
rect 8474 6409 8486 6412
rect 8520 6409 8532 6443
rect 8474 6403 8532 6409
rect 8005 6375 8063 6381
rect 8005 6341 8017 6375
rect 8051 6372 8063 6375
rect 8051 6344 8156 6372
rect 8051 6341 8063 6344
rect 8005 6335 8063 6341
rect 5123 6276 5304 6304
rect 7469 6307 7527 6313
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 7469 6273 7481 6307
rect 7515 6273 7527 6307
rect 7469 6267 7527 6273
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 7834 6304 7840 6316
rect 7699 6276 7840 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 5092 6180 5120 6267
rect 7484 6236 7512 6267
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 8128 6304 8156 6344
rect 8202 6332 8208 6384
rect 8260 6332 8266 6384
rect 8573 6375 8631 6381
rect 8573 6341 8585 6375
rect 8619 6372 8631 6375
rect 8754 6372 8760 6384
rect 8619 6344 8760 6372
rect 8619 6341 8631 6344
rect 8573 6335 8631 6341
rect 8754 6332 8760 6344
rect 8812 6332 8818 6384
rect 8297 6307 8355 6313
rect 8297 6304 8309 6307
rect 8128 6276 8309 6304
rect 8297 6273 8309 6276
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 7484 6208 7880 6236
rect 5074 6128 5080 6180
rect 5132 6128 5138 6180
rect 7852 6177 7880 6208
rect 8312 6180 8340 6267
rect 7837 6171 7895 6177
rect 7837 6137 7849 6171
rect 7883 6168 7895 6171
rect 7926 6168 7932 6180
rect 7883 6140 7932 6168
rect 7883 6137 7895 6140
rect 7837 6131 7895 6137
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 8294 6128 8300 6180
rect 8352 6128 8358 6180
rect 5353 6103 5411 6109
rect 5353 6100 5365 6103
rect 5000 6072 5365 6100
rect 5353 6069 5365 6072
rect 5399 6069 5411 6103
rect 5353 6063 5411 6069
rect 7650 6060 7656 6112
rect 7708 6060 7714 6112
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6100 8079 6103
rect 8202 6100 8208 6112
rect 8067 6072 8208 6100
rect 8067 6069 8079 6072
rect 8021 6063 8079 6069
rect 8202 6060 8208 6072
rect 8260 6100 8266 6112
rect 8404 6100 8432 6267
rect 8260 6072 8432 6100
rect 8260 6060 8266 6072
rect 1104 6010 10120 6032
rect 1104 5958 2077 6010
rect 2129 5958 2141 6010
rect 2193 5958 2205 6010
rect 2257 5958 2269 6010
rect 2321 5958 2333 6010
rect 2385 5958 4331 6010
rect 4383 5958 4395 6010
rect 4447 5958 4459 6010
rect 4511 5958 4523 6010
rect 4575 5958 4587 6010
rect 4639 5958 6585 6010
rect 6637 5958 6649 6010
rect 6701 5958 6713 6010
rect 6765 5958 6777 6010
rect 6829 5958 6841 6010
rect 6893 5958 8839 6010
rect 8891 5958 8903 6010
rect 8955 5958 8967 6010
rect 9019 5958 9031 6010
rect 9083 5958 9095 6010
rect 9147 5958 10120 6010
rect 1104 5936 10120 5958
rect 4706 5856 4712 5908
rect 4764 5856 4770 5908
rect 4801 5899 4859 5905
rect 4801 5865 4813 5899
rect 4847 5896 4859 5899
rect 5074 5896 5080 5908
rect 4847 5868 5080 5896
rect 4847 5865 4859 5868
rect 4801 5859 4859 5865
rect 5074 5856 5080 5868
rect 5132 5856 5138 5908
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8352 5868 9045 5896
rect 8352 5856 8358 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 4724 5760 4752 5856
rect 4890 5788 4896 5840
rect 4948 5788 4954 5840
rect 4172 5732 4752 5760
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 4172 5701 4200 5732
rect 4908 5701 4936 5788
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 5718 5760 5724 5772
rect 5675 5732 5724 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 5718 5720 5724 5732
rect 5776 5720 5782 5772
rect 8570 5720 8576 5772
rect 8628 5760 8634 5772
rect 8628 5732 9168 5760
rect 8628 5720 8634 5732
rect 4157 5695 4215 5701
rect 4157 5692 4169 5695
rect 2746 5664 4169 5692
rect 2746 5624 2774 5664
rect 4157 5661 4169 5664
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5661 4951 5695
rect 4893 5655 4951 5661
rect 1596 5596 2774 5624
rect 1596 5565 1624 5596
rect 4246 5584 4252 5636
rect 4304 5624 4310 5636
rect 4724 5624 4752 5655
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6972 5664 7021 5692
rect 6972 5652 6978 5664
rect 7009 5661 7021 5664
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 8386 5652 8392 5704
rect 8444 5652 8450 5704
rect 8662 5652 8668 5704
rect 8720 5692 8726 5704
rect 9140 5701 9168 5732
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8720 5664 8953 5692
rect 8720 5652 8726 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 4304 5596 4752 5624
rect 7285 5627 7343 5633
rect 4304 5584 4310 5596
rect 7285 5593 7297 5627
rect 7331 5593 7343 5627
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 7285 5587 7343 5593
rect 8772 5596 9413 5624
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5525 1639 5559
rect 1581 5519 1639 5525
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 4065 5559 4123 5565
rect 4065 5556 4077 5559
rect 3936 5528 4077 5556
rect 3936 5516 3942 5528
rect 4065 5525 4077 5528
rect 4111 5556 4123 5559
rect 4890 5556 4896 5568
rect 4111 5528 4896 5556
rect 4111 5525 4123 5528
rect 4065 5519 4123 5525
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 4985 5559 5043 5565
rect 4985 5525 4997 5559
rect 5031 5556 5043 5559
rect 5350 5556 5356 5568
rect 5031 5528 5356 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 7006 5516 7012 5568
rect 7064 5556 7070 5568
rect 7300 5556 7328 5587
rect 8772 5565 8800 5596
rect 9401 5593 9413 5596
rect 9447 5593 9459 5627
rect 9401 5587 9459 5593
rect 7064 5528 7328 5556
rect 8757 5559 8815 5565
rect 7064 5516 7070 5528
rect 8757 5525 8769 5559
rect 8803 5525 8815 5559
rect 8757 5519 8815 5525
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 10042 5556 10048 5568
rect 9723 5528 10048 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 1104 5466 10120 5488
rect 1104 5414 2737 5466
rect 2789 5414 2801 5466
rect 2853 5414 2865 5466
rect 2917 5414 2929 5466
rect 2981 5414 2993 5466
rect 3045 5414 4991 5466
rect 5043 5414 5055 5466
rect 5107 5414 5119 5466
rect 5171 5414 5183 5466
rect 5235 5414 5247 5466
rect 5299 5414 7245 5466
rect 7297 5414 7309 5466
rect 7361 5414 7373 5466
rect 7425 5414 7437 5466
rect 7489 5414 7501 5466
rect 7553 5414 9499 5466
rect 9551 5414 9563 5466
rect 9615 5414 9627 5466
rect 9679 5414 9691 5466
rect 9743 5414 9755 5466
rect 9807 5414 10120 5466
rect 1104 5392 10120 5414
rect 1857 5355 1915 5361
rect 1857 5321 1869 5355
rect 1903 5352 1915 5355
rect 4246 5352 4252 5364
rect 1903 5324 4252 5352
rect 1903 5321 1915 5324
rect 1857 5315 1915 5321
rect 4246 5312 4252 5324
rect 4304 5312 4310 5364
rect 7006 5312 7012 5364
rect 7064 5312 7070 5364
rect 8202 5312 8208 5364
rect 8260 5312 8266 5364
rect 2866 5244 2872 5296
rect 2924 5284 2930 5296
rect 3234 5284 3240 5296
rect 2924 5256 3240 5284
rect 2924 5244 2930 5256
rect 3234 5244 3240 5256
rect 3292 5284 3298 5296
rect 3878 5284 3884 5296
rect 3292 5256 3884 5284
rect 3292 5244 3298 5256
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 4890 5284 4896 5296
rect 4738 5256 4896 5284
rect 4890 5244 4896 5256
rect 4948 5244 4954 5296
rect 5169 5287 5227 5293
rect 5169 5253 5181 5287
rect 5215 5284 5227 5287
rect 8389 5287 8447 5293
rect 5215 5256 6592 5284
rect 5215 5253 5227 5256
rect 5169 5247 5227 5253
rect 3326 5108 3332 5160
rect 3384 5108 3390 5160
rect 3602 5108 3608 5160
rect 3660 5108 3666 5160
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5148 3755 5151
rect 4798 5148 4804 5160
rect 3743 5120 4804 5148
rect 3743 5117 3755 5120
rect 3697 5111 3755 5117
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 5445 5151 5503 5157
rect 5445 5148 5457 5151
rect 5368 5120 5457 5148
rect 3620 5080 3648 5108
rect 3620 5052 4200 5080
rect 4172 5012 4200 5052
rect 5368 5012 5396 5120
rect 5445 5117 5457 5120
rect 5491 5117 5503 5151
rect 5445 5111 5503 5117
rect 6564 5080 6592 5256
rect 6656 5256 7236 5284
rect 6656 5225 6684 5256
rect 7208 5228 7236 5256
rect 7300 5256 7972 5284
rect 7300 5228 7328 5256
rect 7944 5228 7972 5256
rect 8389 5253 8401 5287
rect 8435 5284 8447 5287
rect 8662 5284 8668 5296
rect 8435 5256 8668 5284
rect 8435 5253 8447 5256
rect 8389 5247 8447 5253
rect 8662 5244 8668 5256
rect 8720 5244 8726 5296
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 7190 5176 7196 5228
rect 7248 5176 7254 5228
rect 7282 5176 7288 5228
rect 7340 5176 7346 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 7392 5188 7573 5216
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5148 6975 5151
rect 7098 5148 7104 5160
rect 6963 5120 7104 5148
rect 6963 5117 6975 5120
rect 6917 5111 6975 5117
rect 7098 5108 7104 5120
rect 7156 5148 7162 5160
rect 7392 5148 7420 5188
rect 7561 5185 7573 5188
rect 7607 5216 7619 5219
rect 7607 5188 7788 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7156 5120 7420 5148
rect 7469 5151 7527 5157
rect 7156 5108 7162 5120
rect 7469 5117 7481 5151
rect 7515 5148 7527 5151
rect 7650 5148 7656 5160
rect 7515 5120 7656 5148
rect 7515 5117 7527 5120
rect 7469 5111 7527 5117
rect 7650 5108 7656 5120
rect 7708 5108 7714 5160
rect 7760 5148 7788 5188
rect 7834 5176 7840 5228
rect 7892 5176 7898 5228
rect 7926 5176 7932 5228
rect 7984 5216 7990 5228
rect 8021 5219 8079 5225
rect 8021 5216 8033 5219
rect 7984 5188 8033 5216
rect 7984 5176 7990 5188
rect 8021 5185 8033 5188
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 8570 5176 8576 5228
rect 8628 5176 8634 5228
rect 8113 5151 8171 5157
rect 8113 5148 8125 5151
rect 7760 5120 8125 5148
rect 8113 5117 8125 5120
rect 8159 5117 8171 5151
rect 8113 5111 8171 5117
rect 8662 5080 8668 5092
rect 6564 5052 8668 5080
rect 8662 5040 8668 5052
rect 8720 5040 8726 5092
rect 4172 4984 5396 5012
rect 6454 4972 6460 5024
rect 6512 4972 6518 5024
rect 6825 5015 6883 5021
rect 6825 4981 6837 5015
rect 6871 5012 6883 5015
rect 7282 5012 7288 5024
rect 6871 4984 7288 5012
rect 6871 4981 6883 4984
rect 6825 4975 6883 4981
rect 7282 4972 7288 4984
rect 7340 4972 7346 5024
rect 7650 4972 7656 5024
rect 7708 4972 7714 5024
rect 1104 4922 10120 4944
rect 1104 4870 2077 4922
rect 2129 4870 2141 4922
rect 2193 4870 2205 4922
rect 2257 4870 2269 4922
rect 2321 4870 2333 4922
rect 2385 4870 4331 4922
rect 4383 4870 4395 4922
rect 4447 4870 4459 4922
rect 4511 4870 4523 4922
rect 4575 4870 4587 4922
rect 4639 4870 6585 4922
rect 6637 4870 6649 4922
rect 6701 4870 6713 4922
rect 6765 4870 6777 4922
rect 6829 4870 6841 4922
rect 6893 4870 8839 4922
rect 8891 4870 8903 4922
rect 8955 4870 8967 4922
rect 9019 4870 9031 4922
rect 9083 4870 9095 4922
rect 9147 4870 10120 4922
rect 1104 4848 10120 4870
rect 2406 4768 2412 4820
rect 2464 4808 2470 4820
rect 2866 4808 2872 4820
rect 2464 4780 2872 4808
rect 2464 4768 2470 4780
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 7190 4768 7196 4820
rect 7248 4768 7254 4820
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7834 4808 7840 4820
rect 7607 4780 7840 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7098 4564 7104 4616
rect 7156 4564 7162 4616
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4604 7343 4607
rect 7576 4604 7604 4771
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 7331 4576 7604 4604
rect 7653 4607 7711 4613
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 7742 4604 7748 4616
rect 7699 4576 7748 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 1104 4378 10120 4400
rect 1104 4326 2737 4378
rect 2789 4326 2801 4378
rect 2853 4326 2865 4378
rect 2917 4326 2929 4378
rect 2981 4326 2993 4378
rect 3045 4326 4991 4378
rect 5043 4326 5055 4378
rect 5107 4326 5119 4378
rect 5171 4326 5183 4378
rect 5235 4326 5247 4378
rect 5299 4326 7245 4378
rect 7297 4326 7309 4378
rect 7361 4326 7373 4378
rect 7425 4326 7437 4378
rect 7489 4326 7501 4378
rect 7553 4326 9499 4378
rect 9551 4326 9563 4378
rect 9615 4326 9627 4378
rect 9679 4326 9691 4378
rect 9743 4326 9755 4378
rect 9807 4326 10120 4378
rect 1104 4304 10120 4326
rect 1104 3834 10120 3856
rect 1104 3782 2077 3834
rect 2129 3782 2141 3834
rect 2193 3782 2205 3834
rect 2257 3782 2269 3834
rect 2321 3782 2333 3834
rect 2385 3782 4331 3834
rect 4383 3782 4395 3834
rect 4447 3782 4459 3834
rect 4511 3782 4523 3834
rect 4575 3782 4587 3834
rect 4639 3782 6585 3834
rect 6637 3782 6649 3834
rect 6701 3782 6713 3834
rect 6765 3782 6777 3834
rect 6829 3782 6841 3834
rect 6893 3782 8839 3834
rect 8891 3782 8903 3834
rect 8955 3782 8967 3834
rect 9019 3782 9031 3834
rect 9083 3782 9095 3834
rect 9147 3782 10120 3834
rect 1104 3760 10120 3782
rect 7285 3587 7343 3593
rect 7285 3553 7297 3587
rect 7331 3584 7343 3587
rect 7650 3584 7656 3596
rect 7331 3556 7656 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 7650 3544 7656 3556
rect 7708 3544 7714 3596
rect 6822 3476 6828 3528
rect 6880 3516 6886 3528
rect 7009 3519 7067 3525
rect 7009 3516 7021 3519
rect 6880 3488 7021 3516
rect 6880 3476 6886 3488
rect 7009 3485 7021 3488
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 8754 3340 8760 3392
rect 8812 3340 8818 3392
rect 1104 3290 10120 3312
rect 1104 3238 2737 3290
rect 2789 3238 2801 3290
rect 2853 3238 2865 3290
rect 2917 3238 2929 3290
rect 2981 3238 2993 3290
rect 3045 3238 4991 3290
rect 5043 3238 5055 3290
rect 5107 3238 5119 3290
rect 5171 3238 5183 3290
rect 5235 3238 5247 3290
rect 5299 3238 7245 3290
rect 7297 3238 7309 3290
rect 7361 3238 7373 3290
rect 7425 3238 7437 3290
rect 7489 3238 7501 3290
rect 7553 3238 9499 3290
rect 9551 3238 9563 3290
rect 9615 3238 9627 3290
rect 9679 3238 9691 3290
rect 9743 3238 9755 3290
rect 9807 3238 10120 3290
rect 1104 3216 10120 3238
rect 4890 3136 4896 3188
rect 4948 3176 4954 3188
rect 4948 3148 8432 3176
rect 4948 3136 4954 3148
rect 3694 3068 3700 3120
rect 3752 3068 3758 3120
rect 4908 3108 4936 3136
rect 8404 3120 8432 3148
rect 8570 3136 8576 3188
rect 8628 3136 8634 3188
rect 8754 3136 8760 3188
rect 8812 3136 8818 3188
rect 4830 3080 4936 3108
rect 5261 3111 5319 3117
rect 5261 3077 5273 3111
rect 5307 3108 5319 3111
rect 5350 3108 5356 3120
rect 5307 3080 5356 3108
rect 5307 3077 5319 3080
rect 5261 3071 5319 3077
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 8386 3108 8392 3120
rect 8326 3080 8392 3108
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 1486 3000 1492 3052
rect 1544 3000 1550 3052
rect 8772 3040 8800 3136
rect 9493 3043 9551 3049
rect 9493 3040 9505 3043
rect 8772 3012 9505 3040
rect 9493 3009 9505 3012
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2972 3847 2975
rect 4706 2972 4712 2984
rect 3835 2944 4712 2972
rect 3835 2941 3847 2944
rect 3789 2935 3847 2941
rect 4706 2932 4712 2944
rect 4764 2932 4770 2984
rect 5537 2975 5595 2981
rect 5537 2941 5549 2975
rect 5583 2972 5595 2975
rect 6822 2972 6828 2984
rect 5583 2944 6828 2972
rect 5583 2941 5595 2944
rect 5537 2935 5595 2941
rect 3602 2904 3608 2916
rect 2884 2876 3608 2904
rect 2884 2848 2912 2876
rect 3602 2864 3608 2876
rect 3660 2904 3666 2916
rect 3660 2876 4108 2904
rect 3660 2864 3666 2876
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 992 2808 1593 2836
rect 992 2796 998 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 2409 2839 2467 2845
rect 2409 2805 2421 2839
rect 2455 2836 2467 2839
rect 2866 2836 2872 2848
rect 2455 2808 2872 2836
rect 2455 2805 2467 2808
rect 2409 2799 2467 2805
rect 2866 2796 2872 2808
rect 2924 2796 2930 2848
rect 4080 2836 4108 2876
rect 5552 2836 5580 2935
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 7101 2975 7159 2981
rect 7101 2941 7113 2975
rect 7147 2972 7159 2975
rect 8478 2972 8484 2984
rect 7147 2944 8484 2972
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 4080 2808 5580 2836
rect 9674 2796 9680 2848
rect 9732 2796 9738 2848
rect 1104 2746 10120 2768
rect 1104 2694 2077 2746
rect 2129 2694 2141 2746
rect 2193 2694 2205 2746
rect 2257 2694 2269 2746
rect 2321 2694 2333 2746
rect 2385 2694 4331 2746
rect 4383 2694 4395 2746
rect 4447 2694 4459 2746
rect 4511 2694 4523 2746
rect 4575 2694 4587 2746
rect 4639 2694 6585 2746
rect 6637 2694 6649 2746
rect 6701 2694 6713 2746
rect 6765 2694 6777 2746
rect 6829 2694 6841 2746
rect 6893 2694 8839 2746
rect 8891 2694 8903 2746
rect 8955 2694 8967 2746
rect 9019 2694 9031 2746
rect 9083 2694 9095 2746
rect 9147 2694 10120 2746
rect 1104 2672 10120 2694
rect 1397 2635 1455 2641
rect 1397 2601 1409 2635
rect 1443 2632 1455 2635
rect 1486 2632 1492 2644
rect 1443 2604 1492 2632
rect 1443 2601 1455 2604
rect 1397 2595 1455 2601
rect 1486 2592 1492 2604
rect 1544 2592 1550 2644
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 3326 2632 3332 2644
rect 3283 2604 3332 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 6454 2592 6460 2644
rect 6512 2592 6518 2644
rect 8478 2592 8484 2644
rect 8536 2592 8542 2644
rect 8662 2592 8668 2644
rect 8720 2632 8726 2644
rect 9585 2635 9643 2641
rect 9585 2632 9597 2635
rect 8720 2604 9597 2632
rect 8720 2592 8726 2604
rect 9585 2601 9597 2604
rect 9631 2601 9643 2635
rect 9585 2595 9643 2601
rect 2866 2456 2872 2508
rect 2924 2496 2930 2508
rect 3145 2499 3203 2505
rect 3145 2496 3157 2499
rect 2924 2468 3157 2496
rect 2924 2456 2930 2468
rect 3145 2465 3157 2468
rect 3191 2465 3203 2499
rect 6472 2496 6500 2592
rect 3145 2459 3203 2465
rect 3344 2468 6500 2496
rect 2406 2320 2412 2372
rect 2464 2320 2470 2372
rect 2869 2363 2927 2369
rect 2869 2329 2881 2363
rect 2915 2360 2927 2363
rect 3344 2360 3372 2468
rect 3421 2431 3479 2437
rect 3421 2397 3433 2431
rect 3467 2397 3479 2431
rect 3421 2391 3479 2397
rect 2915 2332 3372 2360
rect 2915 2329 2927 2332
rect 2869 2323 2927 2329
rect 14 2252 20 2304
rect 72 2292 78 2304
rect 3436 2292 3464 2391
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 5169 2431 5227 2437
rect 5169 2428 5181 2431
rect 4764 2400 5181 2428
rect 4764 2388 4770 2400
rect 5169 2397 5181 2400
rect 5215 2397 5227 2431
rect 5169 2391 5227 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 8444 2400 8677 2428
rect 8444 2388 8450 2400
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 9769 2431 9827 2437
rect 9769 2397 9781 2431
rect 9815 2428 9827 2431
rect 10962 2428 10968 2440
rect 9815 2400 10968 2428
rect 9815 2397 9827 2400
rect 9769 2391 9827 2397
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 72 2264 3464 2292
rect 5261 2295 5319 2301
rect 72 2252 78 2264
rect 5261 2261 5273 2295
rect 5307 2292 5319 2295
rect 5350 2292 5356 2304
rect 5307 2264 5356 2292
rect 5307 2261 5319 2264
rect 5261 2255 5319 2261
rect 5350 2252 5356 2264
rect 5408 2252 5414 2304
rect 1104 2202 10120 2224
rect 1104 2150 2737 2202
rect 2789 2150 2801 2202
rect 2853 2150 2865 2202
rect 2917 2150 2929 2202
rect 2981 2150 2993 2202
rect 3045 2150 4991 2202
rect 5043 2150 5055 2202
rect 5107 2150 5119 2202
rect 5171 2150 5183 2202
rect 5235 2150 5247 2202
rect 5299 2150 7245 2202
rect 7297 2150 7309 2202
rect 7361 2150 7373 2202
rect 7425 2150 7437 2202
rect 7489 2150 7501 2202
rect 7553 2150 9499 2202
rect 9551 2150 9563 2202
rect 9615 2150 9627 2202
rect 9679 2150 9691 2202
rect 9743 2150 9755 2202
rect 9807 2150 10120 2202
rect 1104 2128 10120 2150
<< via1 >>
rect 2737 10854 2789 10906
rect 2801 10854 2853 10906
rect 2865 10854 2917 10906
rect 2929 10854 2981 10906
rect 2993 10854 3045 10906
rect 4991 10854 5043 10906
rect 5055 10854 5107 10906
rect 5119 10854 5171 10906
rect 5183 10854 5235 10906
rect 5247 10854 5299 10906
rect 7245 10854 7297 10906
rect 7309 10854 7361 10906
rect 7373 10854 7425 10906
rect 7437 10854 7489 10906
rect 7501 10854 7553 10906
rect 9499 10854 9551 10906
rect 9563 10854 9615 10906
rect 9627 10854 9679 10906
rect 9691 10854 9743 10906
rect 9755 10854 9807 10906
rect 1308 10752 1360 10804
rect 7104 10752 7156 10804
rect 9312 10752 9364 10804
rect 9864 10752 9916 10804
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 1952 10659 2004 10668
rect 1952 10625 1961 10659
rect 1961 10625 1995 10659
rect 1995 10625 2004 10659
rect 1952 10616 2004 10625
rect 3884 10616 3936 10668
rect 3608 10548 3660 10600
rect 5264 10659 5316 10668
rect 5264 10625 5273 10659
rect 5273 10625 5307 10659
rect 5307 10625 5316 10659
rect 5264 10616 5316 10625
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 5816 10616 5868 10668
rect 1952 10412 2004 10464
rect 3976 10455 4028 10464
rect 3976 10421 3985 10455
rect 3985 10421 4019 10455
rect 4019 10421 4028 10455
rect 3976 10412 4028 10421
rect 4252 10412 4304 10464
rect 5540 10412 5592 10464
rect 5632 10412 5684 10464
rect 6368 10412 6420 10464
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 9588 10455 9640 10464
rect 9588 10421 9597 10455
rect 9597 10421 9631 10455
rect 9631 10421 9640 10455
rect 9588 10412 9640 10421
rect 2077 10310 2129 10362
rect 2141 10310 2193 10362
rect 2205 10310 2257 10362
rect 2269 10310 2321 10362
rect 2333 10310 2385 10362
rect 4331 10310 4383 10362
rect 4395 10310 4447 10362
rect 4459 10310 4511 10362
rect 4523 10310 4575 10362
rect 4587 10310 4639 10362
rect 6585 10310 6637 10362
rect 6649 10310 6701 10362
rect 6713 10310 6765 10362
rect 6777 10310 6829 10362
rect 6841 10310 6893 10362
rect 8839 10310 8891 10362
rect 8903 10310 8955 10362
rect 8967 10310 9019 10362
rect 9031 10310 9083 10362
rect 9095 10310 9147 10362
rect 1952 10208 2004 10260
rect 3608 10251 3660 10260
rect 3608 10217 3617 10251
rect 3617 10217 3651 10251
rect 3651 10217 3660 10251
rect 3608 10208 3660 10217
rect 5264 10208 5316 10260
rect 9312 10208 9364 10260
rect 9588 10208 9640 10260
rect 3424 10072 3476 10124
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 4528 10004 4580 10013
rect 5172 10072 5224 10124
rect 5264 10072 5316 10124
rect 6460 10072 6512 10124
rect 4712 9936 4764 9988
rect 7104 9936 7156 9988
rect 4160 9911 4212 9920
rect 4160 9877 4169 9911
rect 4169 9877 4203 9911
rect 4203 9877 4212 9911
rect 4160 9868 4212 9877
rect 5632 9868 5684 9920
rect 8668 9911 8720 9920
rect 8668 9877 8677 9911
rect 8677 9877 8711 9911
rect 8711 9877 8720 9911
rect 8668 9868 8720 9877
rect 2737 9766 2789 9818
rect 2801 9766 2853 9818
rect 2865 9766 2917 9818
rect 2929 9766 2981 9818
rect 2993 9766 3045 9818
rect 4991 9766 5043 9818
rect 5055 9766 5107 9818
rect 5119 9766 5171 9818
rect 5183 9766 5235 9818
rect 5247 9766 5299 9818
rect 7245 9766 7297 9818
rect 7309 9766 7361 9818
rect 7373 9766 7425 9818
rect 7437 9766 7489 9818
rect 7501 9766 7553 9818
rect 9499 9766 9551 9818
rect 9563 9766 9615 9818
rect 9627 9766 9679 9818
rect 9691 9766 9743 9818
rect 9755 9766 9807 9818
rect 1492 9664 1544 9716
rect 4252 9664 4304 9716
rect 4160 9596 4212 9648
rect 4528 9664 4580 9716
rect 5632 9707 5684 9716
rect 5632 9673 5659 9707
rect 5659 9673 5684 9707
rect 5632 9664 5684 9673
rect 5816 9639 5868 9648
rect 5816 9605 5825 9639
rect 5825 9605 5859 9639
rect 5859 9605 5868 9639
rect 5816 9596 5868 9605
rect 3424 9460 3476 9512
rect 4436 9460 4488 9512
rect 3240 9324 3292 9376
rect 4804 9367 4856 9376
rect 4804 9333 4813 9367
rect 4813 9333 4847 9367
rect 4847 9333 4856 9367
rect 4804 9324 4856 9333
rect 5172 9324 5224 9376
rect 5540 9324 5592 9376
rect 2077 9222 2129 9274
rect 2141 9222 2193 9274
rect 2205 9222 2257 9274
rect 2269 9222 2321 9274
rect 2333 9222 2385 9274
rect 4331 9222 4383 9274
rect 4395 9222 4447 9274
rect 4459 9222 4511 9274
rect 4523 9222 4575 9274
rect 4587 9222 4639 9274
rect 6585 9222 6637 9274
rect 6649 9222 6701 9274
rect 6713 9222 6765 9274
rect 6777 9222 6829 9274
rect 6841 9222 6893 9274
rect 8839 9222 8891 9274
rect 8903 9222 8955 9274
rect 8967 9222 9019 9274
rect 9031 9222 9083 9274
rect 9095 9222 9147 9274
rect 4804 9120 4856 9172
rect 6920 9120 6972 9172
rect 6644 8916 6696 8968
rect 10140 8916 10192 8968
rect 1492 8891 1544 8900
rect 1492 8857 1501 8891
rect 1501 8857 1535 8891
rect 1535 8857 1544 8891
rect 1492 8848 1544 8857
rect 940 8780 992 8832
rect 6276 8780 6328 8832
rect 8852 8780 8904 8832
rect 2737 8678 2789 8730
rect 2801 8678 2853 8730
rect 2865 8678 2917 8730
rect 2929 8678 2981 8730
rect 2993 8678 3045 8730
rect 4991 8678 5043 8730
rect 5055 8678 5107 8730
rect 5119 8678 5171 8730
rect 5183 8678 5235 8730
rect 5247 8678 5299 8730
rect 7245 8678 7297 8730
rect 7309 8678 7361 8730
rect 7373 8678 7425 8730
rect 7437 8678 7489 8730
rect 7501 8678 7553 8730
rect 9499 8678 9551 8730
rect 9563 8678 9615 8730
rect 9627 8678 9679 8730
rect 9691 8678 9743 8730
rect 9755 8678 9807 8730
rect 1492 8576 1544 8628
rect 4712 8576 4764 8628
rect 3240 8508 3292 8560
rect 3976 8508 4028 8560
rect 7104 8576 7156 8628
rect 8208 8576 8260 8628
rect 8852 8576 8904 8628
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 4160 8372 4212 8424
rect 4712 8372 4764 8424
rect 8392 8415 8444 8424
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 6644 8347 6696 8356
rect 6644 8313 6653 8347
rect 6653 8313 6687 8347
rect 6687 8313 6696 8347
rect 6644 8304 6696 8313
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 5908 8236 5960 8288
rect 2077 8134 2129 8186
rect 2141 8134 2193 8186
rect 2205 8134 2257 8186
rect 2269 8134 2321 8186
rect 2333 8134 2385 8186
rect 4331 8134 4383 8186
rect 4395 8134 4447 8186
rect 4459 8134 4511 8186
rect 4523 8134 4575 8186
rect 4587 8134 4639 8186
rect 6585 8134 6637 8186
rect 6649 8134 6701 8186
rect 6713 8134 6765 8186
rect 6777 8134 6829 8186
rect 6841 8134 6893 8186
rect 8839 8134 8891 8186
rect 8903 8134 8955 8186
rect 8967 8134 9019 8186
rect 9031 8134 9083 8186
rect 9095 8134 9147 8186
rect 3424 8032 3476 8084
rect 6460 8032 6512 8084
rect 5172 7896 5224 7948
rect 5724 7939 5776 7948
rect 5724 7905 5733 7939
rect 5733 7905 5767 7939
rect 5767 7905 5776 7939
rect 5724 7896 5776 7905
rect 8392 8032 8444 8084
rect 5908 7828 5960 7880
rect 6276 7828 6328 7880
rect 4252 7760 4304 7812
rect 5448 7760 5500 7812
rect 6368 7760 6420 7812
rect 7104 7760 7156 7812
rect 4896 7735 4948 7744
rect 4896 7701 4905 7735
rect 4905 7701 4939 7735
rect 4939 7701 4948 7735
rect 4896 7692 4948 7701
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 2737 7590 2789 7642
rect 2801 7590 2853 7642
rect 2865 7590 2917 7642
rect 2929 7590 2981 7642
rect 2993 7590 3045 7642
rect 4991 7590 5043 7642
rect 5055 7590 5107 7642
rect 5119 7590 5171 7642
rect 5183 7590 5235 7642
rect 5247 7590 5299 7642
rect 7245 7590 7297 7642
rect 7309 7590 7361 7642
rect 7373 7590 7425 7642
rect 7437 7590 7489 7642
rect 7501 7590 7553 7642
rect 9499 7590 9551 7642
rect 9563 7590 9615 7642
rect 9627 7590 9679 7642
rect 9691 7590 9743 7642
rect 9755 7590 9807 7642
rect 3424 7488 3476 7540
rect 4160 7488 4212 7540
rect 4896 7488 4948 7540
rect 5356 7488 5408 7540
rect 4160 7352 4212 7404
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 5540 7352 5592 7404
rect 8300 7352 8352 7404
rect 4896 7148 4948 7200
rect 8760 7148 8812 7200
rect 2077 7046 2129 7098
rect 2141 7046 2193 7098
rect 2205 7046 2257 7098
rect 2269 7046 2321 7098
rect 2333 7046 2385 7098
rect 4331 7046 4383 7098
rect 4395 7046 4447 7098
rect 4459 7046 4511 7098
rect 4523 7046 4575 7098
rect 4587 7046 4639 7098
rect 6585 7046 6637 7098
rect 6649 7046 6701 7098
rect 6713 7046 6765 7098
rect 6777 7046 6829 7098
rect 6841 7046 6893 7098
rect 8839 7046 8891 7098
rect 8903 7046 8955 7098
rect 8967 7046 9019 7098
rect 9031 7046 9083 7098
rect 9095 7046 9147 7098
rect 4160 6944 4212 6996
rect 5540 6944 5592 6996
rect 4804 6808 4856 6860
rect 4896 6740 4948 6792
rect 4160 6672 4212 6724
rect 2737 6502 2789 6554
rect 2801 6502 2853 6554
rect 2865 6502 2917 6554
rect 2929 6502 2981 6554
rect 2993 6502 3045 6554
rect 4991 6502 5043 6554
rect 5055 6502 5107 6554
rect 5119 6502 5171 6554
rect 5183 6502 5235 6554
rect 5247 6502 5299 6554
rect 7245 6502 7297 6554
rect 7309 6502 7361 6554
rect 7373 6502 7425 6554
rect 7437 6502 7489 6554
rect 7501 6502 7553 6554
rect 9499 6502 9551 6554
rect 9563 6502 9615 6554
rect 9627 6502 9679 6554
rect 9691 6502 9743 6554
rect 9755 6502 9807 6554
rect 4252 6400 4304 6452
rect 4896 6400 4948 6452
rect 5080 6400 5132 6452
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 4252 6264 4304 6316
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 4804 6264 4856 6273
rect 4896 6196 4948 6248
rect 7840 6264 7892 6316
rect 8208 6375 8260 6384
rect 8208 6341 8217 6375
rect 8217 6341 8251 6375
rect 8251 6341 8260 6375
rect 8208 6332 8260 6341
rect 8760 6332 8812 6384
rect 5080 6128 5132 6180
rect 7932 6128 7984 6180
rect 8300 6128 8352 6180
rect 7656 6103 7708 6112
rect 7656 6069 7665 6103
rect 7665 6069 7699 6103
rect 7699 6069 7708 6103
rect 7656 6060 7708 6069
rect 8208 6060 8260 6112
rect 2077 5958 2129 6010
rect 2141 5958 2193 6010
rect 2205 5958 2257 6010
rect 2269 5958 2321 6010
rect 2333 5958 2385 6010
rect 4331 5958 4383 6010
rect 4395 5958 4447 6010
rect 4459 5958 4511 6010
rect 4523 5958 4575 6010
rect 4587 5958 4639 6010
rect 6585 5958 6637 6010
rect 6649 5958 6701 6010
rect 6713 5958 6765 6010
rect 6777 5958 6829 6010
rect 6841 5958 6893 6010
rect 8839 5958 8891 6010
rect 8903 5958 8955 6010
rect 8967 5958 9019 6010
rect 9031 5958 9083 6010
rect 9095 5958 9147 6010
rect 4712 5856 4764 5908
rect 5080 5856 5132 5908
rect 8300 5856 8352 5908
rect 4896 5788 4948 5840
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 5724 5720 5776 5772
rect 8576 5720 8628 5772
rect 4252 5584 4304 5636
rect 6920 5652 6972 5704
rect 8392 5652 8444 5704
rect 8668 5652 8720 5704
rect 3884 5516 3936 5568
rect 4896 5516 4948 5568
rect 5356 5516 5408 5568
rect 7012 5516 7064 5568
rect 10048 5516 10100 5568
rect 2737 5414 2789 5466
rect 2801 5414 2853 5466
rect 2865 5414 2917 5466
rect 2929 5414 2981 5466
rect 2993 5414 3045 5466
rect 4991 5414 5043 5466
rect 5055 5414 5107 5466
rect 5119 5414 5171 5466
rect 5183 5414 5235 5466
rect 5247 5414 5299 5466
rect 7245 5414 7297 5466
rect 7309 5414 7361 5466
rect 7373 5414 7425 5466
rect 7437 5414 7489 5466
rect 7501 5414 7553 5466
rect 9499 5414 9551 5466
rect 9563 5414 9615 5466
rect 9627 5414 9679 5466
rect 9691 5414 9743 5466
rect 9755 5414 9807 5466
rect 4252 5312 4304 5364
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 8208 5355 8260 5364
rect 8208 5321 8217 5355
rect 8217 5321 8251 5355
rect 8251 5321 8260 5355
rect 8208 5312 8260 5321
rect 2872 5244 2924 5296
rect 3240 5244 3292 5296
rect 3884 5244 3936 5296
rect 4896 5244 4948 5296
rect 3332 5151 3384 5160
rect 3332 5117 3341 5151
rect 3341 5117 3375 5151
rect 3375 5117 3384 5151
rect 3332 5108 3384 5117
rect 3608 5151 3660 5160
rect 3608 5117 3617 5151
rect 3617 5117 3651 5151
rect 3651 5117 3660 5151
rect 3608 5108 3660 5117
rect 4804 5108 4856 5160
rect 8668 5244 8720 5296
rect 7196 5219 7248 5228
rect 7196 5185 7205 5219
rect 7205 5185 7239 5219
rect 7239 5185 7248 5219
rect 7196 5176 7248 5185
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 7104 5108 7156 5160
rect 7656 5108 7708 5160
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 7932 5176 7984 5228
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 8668 5040 8720 5092
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 7288 4972 7340 5024
rect 7656 5015 7708 5024
rect 7656 4981 7665 5015
rect 7665 4981 7699 5015
rect 7699 4981 7708 5015
rect 7656 4972 7708 4981
rect 2077 4870 2129 4922
rect 2141 4870 2193 4922
rect 2205 4870 2257 4922
rect 2269 4870 2321 4922
rect 2333 4870 2385 4922
rect 4331 4870 4383 4922
rect 4395 4870 4447 4922
rect 4459 4870 4511 4922
rect 4523 4870 4575 4922
rect 4587 4870 4639 4922
rect 6585 4870 6637 4922
rect 6649 4870 6701 4922
rect 6713 4870 6765 4922
rect 6777 4870 6829 4922
rect 6841 4870 6893 4922
rect 8839 4870 8891 4922
rect 8903 4870 8955 4922
rect 8967 4870 9019 4922
rect 9031 4870 9083 4922
rect 9095 4870 9147 4922
rect 2412 4768 2464 4820
rect 2872 4768 2924 4820
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 7104 4607 7156 4616
rect 7104 4573 7113 4607
rect 7113 4573 7147 4607
rect 7147 4573 7156 4607
rect 7104 4564 7156 4573
rect 7840 4768 7892 4820
rect 7748 4564 7800 4616
rect 2737 4326 2789 4378
rect 2801 4326 2853 4378
rect 2865 4326 2917 4378
rect 2929 4326 2981 4378
rect 2993 4326 3045 4378
rect 4991 4326 5043 4378
rect 5055 4326 5107 4378
rect 5119 4326 5171 4378
rect 5183 4326 5235 4378
rect 5247 4326 5299 4378
rect 7245 4326 7297 4378
rect 7309 4326 7361 4378
rect 7373 4326 7425 4378
rect 7437 4326 7489 4378
rect 7501 4326 7553 4378
rect 9499 4326 9551 4378
rect 9563 4326 9615 4378
rect 9627 4326 9679 4378
rect 9691 4326 9743 4378
rect 9755 4326 9807 4378
rect 2077 3782 2129 3834
rect 2141 3782 2193 3834
rect 2205 3782 2257 3834
rect 2269 3782 2321 3834
rect 2333 3782 2385 3834
rect 4331 3782 4383 3834
rect 4395 3782 4447 3834
rect 4459 3782 4511 3834
rect 4523 3782 4575 3834
rect 4587 3782 4639 3834
rect 6585 3782 6637 3834
rect 6649 3782 6701 3834
rect 6713 3782 6765 3834
rect 6777 3782 6829 3834
rect 6841 3782 6893 3834
rect 8839 3782 8891 3834
rect 8903 3782 8955 3834
rect 8967 3782 9019 3834
rect 9031 3782 9083 3834
rect 9095 3782 9147 3834
rect 7656 3544 7708 3596
rect 6828 3476 6880 3528
rect 8392 3476 8444 3528
rect 8760 3383 8812 3392
rect 8760 3349 8769 3383
rect 8769 3349 8803 3383
rect 8803 3349 8812 3383
rect 8760 3340 8812 3349
rect 2737 3238 2789 3290
rect 2801 3238 2853 3290
rect 2865 3238 2917 3290
rect 2929 3238 2981 3290
rect 2993 3238 3045 3290
rect 4991 3238 5043 3290
rect 5055 3238 5107 3290
rect 5119 3238 5171 3290
rect 5183 3238 5235 3290
rect 5247 3238 5299 3290
rect 7245 3238 7297 3290
rect 7309 3238 7361 3290
rect 7373 3238 7425 3290
rect 7437 3238 7489 3290
rect 7501 3238 7553 3290
rect 9499 3238 9551 3290
rect 9563 3238 9615 3290
rect 9627 3238 9679 3290
rect 9691 3238 9743 3290
rect 9755 3238 9807 3290
rect 4896 3136 4948 3188
rect 3700 3111 3752 3120
rect 3700 3077 3709 3111
rect 3709 3077 3743 3111
rect 3743 3077 3752 3111
rect 3700 3068 3752 3077
rect 8576 3179 8628 3188
rect 8576 3145 8585 3179
rect 8585 3145 8619 3179
rect 8619 3145 8628 3179
rect 8576 3136 8628 3145
rect 8760 3136 8812 3188
rect 5356 3068 5408 3120
rect 8392 3068 8444 3120
rect 1492 3043 1544 3052
rect 1492 3009 1501 3043
rect 1501 3009 1535 3043
rect 1535 3009 1544 3043
rect 1492 3000 1544 3009
rect 4712 2932 4764 2984
rect 6828 2975 6880 2984
rect 3608 2864 3660 2916
rect 940 2796 992 2848
rect 2872 2796 2924 2848
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 8484 2932 8536 2984
rect 9680 2839 9732 2848
rect 9680 2805 9689 2839
rect 9689 2805 9723 2839
rect 9723 2805 9732 2839
rect 9680 2796 9732 2805
rect 2077 2694 2129 2746
rect 2141 2694 2193 2746
rect 2205 2694 2257 2746
rect 2269 2694 2321 2746
rect 2333 2694 2385 2746
rect 4331 2694 4383 2746
rect 4395 2694 4447 2746
rect 4459 2694 4511 2746
rect 4523 2694 4575 2746
rect 4587 2694 4639 2746
rect 6585 2694 6637 2746
rect 6649 2694 6701 2746
rect 6713 2694 6765 2746
rect 6777 2694 6829 2746
rect 6841 2694 6893 2746
rect 8839 2694 8891 2746
rect 8903 2694 8955 2746
rect 8967 2694 9019 2746
rect 9031 2694 9083 2746
rect 9095 2694 9147 2746
rect 1492 2592 1544 2644
rect 3332 2592 3384 2644
rect 6460 2592 6512 2644
rect 8484 2635 8536 2644
rect 8484 2601 8493 2635
rect 8493 2601 8527 2635
rect 8527 2601 8536 2635
rect 8484 2592 8536 2601
rect 8668 2592 8720 2644
rect 2872 2456 2924 2508
rect 2412 2320 2464 2372
rect 20 2252 72 2304
rect 4712 2388 4764 2440
rect 8392 2388 8444 2440
rect 10968 2388 11020 2440
rect 5356 2252 5408 2304
rect 2737 2150 2789 2202
rect 2801 2150 2853 2202
rect 2865 2150 2917 2202
rect 2929 2150 2981 2202
rect 2993 2150 3045 2202
rect 4991 2150 5043 2202
rect 5055 2150 5107 2202
rect 5119 2150 5171 2202
rect 5183 2150 5235 2202
rect 5247 2150 5299 2202
rect 7245 2150 7297 2202
rect 7309 2150 7361 2202
rect 7373 2150 7425 2202
rect 7437 2150 7489 2202
rect 7501 2150 7553 2202
rect 9499 2150 9551 2202
rect 9563 2150 9615 2202
rect 9627 2150 9679 2202
rect 9691 2150 9743 2202
rect 9755 2150 9807 2202
<< metal2 >>
rect 1306 12639 1362 13439
rect 3882 12639 3938 13439
rect 7102 12639 7158 13439
rect 9678 12639 9734 13439
rect 1320 10810 1348 12639
rect 1950 11656 2006 11665
rect 1950 11591 2006 11600
rect 1308 10804 1360 10810
rect 1308 10746 1360 10752
rect 1964 10674 1992 11591
rect 2737 10908 3045 10917
rect 2737 10906 2743 10908
rect 2799 10906 2823 10908
rect 2879 10906 2903 10908
rect 2959 10906 2983 10908
rect 3039 10906 3045 10908
rect 2799 10854 2801 10906
rect 2981 10854 2983 10906
rect 2737 10852 2743 10854
rect 2799 10852 2823 10854
rect 2879 10852 2903 10854
rect 2959 10852 2983 10854
rect 3039 10852 3045 10854
rect 2737 10843 3045 10852
rect 3896 10674 3924 12639
rect 4991 10908 5299 10917
rect 4991 10906 4997 10908
rect 5053 10906 5077 10908
rect 5133 10906 5157 10908
rect 5213 10906 5237 10908
rect 5293 10906 5299 10908
rect 5053 10854 5055 10906
rect 5235 10854 5237 10906
rect 4991 10852 4997 10854
rect 5053 10852 5077 10854
rect 5133 10852 5157 10854
rect 5213 10852 5237 10854
rect 5293 10852 5299 10854
rect 4991 10843 5299 10852
rect 7116 10810 7144 12639
rect 9310 11656 9366 11665
rect 9692 11642 9720 12639
rect 9692 11614 9904 11642
rect 9310 11591 9366 11600
rect 7245 10908 7553 10917
rect 7245 10906 7251 10908
rect 7307 10906 7331 10908
rect 7387 10906 7411 10908
rect 7467 10906 7491 10908
rect 7547 10906 7553 10908
rect 7307 10854 7309 10906
rect 7489 10854 7491 10906
rect 7245 10852 7251 10854
rect 7307 10852 7331 10854
rect 7387 10852 7411 10854
rect 7467 10852 7491 10854
rect 7547 10852 7553 10854
rect 7245 10843 7553 10852
rect 9324 10810 9352 11591
rect 9499 10908 9807 10917
rect 9499 10906 9505 10908
rect 9561 10906 9585 10908
rect 9641 10906 9665 10908
rect 9721 10906 9745 10908
rect 9801 10906 9807 10908
rect 9561 10854 9563 10906
rect 9743 10854 9745 10906
rect 9499 10852 9505 10854
rect 9561 10852 9585 10854
rect 9641 10852 9665 10854
rect 9721 10852 9745 10854
rect 9801 10852 9807 10854
rect 9499 10843 9807 10852
rect 9876 10810 9904 11614
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9864 10804 9916 10810
rect 9864 10746 9916 10752
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 1504 9722 1532 10610
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 10266 1992 10406
rect 2077 10364 2385 10373
rect 2077 10362 2083 10364
rect 2139 10362 2163 10364
rect 2219 10362 2243 10364
rect 2299 10362 2323 10364
rect 2379 10362 2385 10364
rect 2139 10310 2141 10362
rect 2321 10310 2323 10362
rect 2077 10308 2083 10310
rect 2139 10308 2163 10310
rect 2219 10308 2243 10310
rect 2299 10308 2323 10310
rect 2379 10308 2385 10310
rect 2077 10299 2385 10308
rect 3620 10266 3648 10542
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 2737 9820 3045 9829
rect 2737 9818 2743 9820
rect 2799 9818 2823 9820
rect 2879 9818 2903 9820
rect 2959 9818 2983 9820
rect 3039 9818 3045 9820
rect 2799 9766 2801 9818
rect 2981 9766 2983 9818
rect 2737 9764 2743 9766
rect 2799 9764 2823 9766
rect 2879 9764 2903 9766
rect 2959 9764 2983 9766
rect 3039 9764 3045 9766
rect 2737 9755 3045 9764
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 3436 9518 3464 10066
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 2077 9276 2385 9285
rect 2077 9274 2083 9276
rect 2139 9274 2163 9276
rect 2219 9274 2243 9276
rect 2299 9274 2323 9276
rect 2379 9274 2385 9276
rect 2139 9222 2141 9274
rect 2321 9222 2323 9274
rect 2077 9220 2083 9222
rect 2139 9220 2163 9222
rect 2219 9220 2243 9222
rect 2299 9220 2323 9222
rect 2379 9220 2385 9222
rect 2077 9211 2385 9220
rect 938 8936 994 8945
rect 938 8871 994 8880
rect 1492 8900 1544 8906
rect 952 8838 980 8871
rect 1492 8842 1544 8848
rect 940 8832 992 8838
rect 940 8774 992 8780
rect 1504 8634 1532 8842
rect 2737 8732 3045 8741
rect 2737 8730 2743 8732
rect 2799 8730 2823 8732
rect 2879 8730 2903 8732
rect 2959 8730 2983 8732
rect 3039 8730 3045 8732
rect 2799 8678 2801 8730
rect 2981 8678 2983 8730
rect 2737 8676 2743 8678
rect 2799 8676 2823 8678
rect 2879 8676 2903 8678
rect 2959 8676 2983 8678
rect 3039 8676 3045 8678
rect 2737 8667 3045 8676
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 3252 8566 3280 9318
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 2077 8188 2385 8197
rect 2077 8186 2083 8188
rect 2139 8186 2163 8188
rect 2219 8186 2243 8188
rect 2299 8186 2323 8188
rect 2379 8186 2385 8188
rect 2139 8134 2141 8186
rect 2321 8134 2323 8186
rect 2077 8132 2083 8134
rect 2139 8132 2163 8134
rect 2219 8132 2243 8134
rect 2299 8132 2323 8134
rect 2379 8132 2385 8134
rect 2077 8123 2385 8132
rect 2737 7644 3045 7653
rect 2737 7642 2743 7644
rect 2799 7642 2823 7644
rect 2879 7642 2903 7644
rect 2959 7642 2983 7644
rect 3039 7642 3045 7644
rect 2799 7590 2801 7642
rect 2981 7590 2983 7642
rect 2737 7588 2743 7590
rect 2799 7588 2823 7590
rect 2879 7588 2903 7590
rect 2959 7588 2983 7590
rect 3039 7588 3045 7590
rect 2737 7579 3045 7588
rect 2077 7100 2385 7109
rect 2077 7098 2083 7100
rect 2139 7098 2163 7100
rect 2219 7098 2243 7100
rect 2299 7098 2323 7100
rect 2379 7098 2385 7100
rect 2139 7046 2141 7098
rect 2321 7046 2323 7098
rect 2077 7044 2083 7046
rect 2139 7044 2163 7046
rect 2219 7044 2243 7046
rect 2299 7044 2323 7046
rect 2379 7044 2385 7046
rect 2077 7035 2385 7044
rect 2737 6556 3045 6565
rect 2737 6554 2743 6556
rect 2799 6554 2823 6556
rect 2879 6554 2903 6556
rect 2959 6554 2983 6556
rect 3039 6554 3045 6556
rect 2799 6502 2801 6554
rect 2981 6502 2983 6554
rect 2737 6500 2743 6502
rect 2799 6500 2823 6502
rect 2879 6500 2903 6502
rect 2959 6500 2983 6502
rect 3039 6500 3045 6502
rect 2737 6491 3045 6500
rect 2077 6012 2385 6021
rect 2077 6010 2083 6012
rect 2139 6010 2163 6012
rect 2219 6010 2243 6012
rect 2299 6010 2323 6012
rect 2379 6010 2385 6012
rect 2139 5958 2141 6010
rect 2321 5958 2323 6010
rect 2077 5956 2083 5958
rect 2139 5956 2163 5958
rect 2219 5956 2243 5958
rect 2299 5956 2323 5958
rect 2379 5956 2385 5958
rect 2077 5947 2385 5956
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 2737 5468 3045 5477
rect 2737 5466 2743 5468
rect 2799 5466 2823 5468
rect 2879 5466 2903 5468
rect 2959 5466 2983 5468
rect 3039 5466 3045 5468
rect 2799 5414 2801 5466
rect 2981 5414 2983 5466
rect 2737 5412 2743 5414
rect 2799 5412 2823 5414
rect 2879 5412 2903 5414
rect 2959 5412 2983 5414
rect 3039 5412 3045 5414
rect 2737 5403 3045 5412
rect 3252 5302 3280 8502
rect 3436 8430 3464 9454
rect 3988 8566 4016 10406
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4172 9654 4200 9862
rect 4264 9722 4292 10406
rect 4331 10364 4639 10373
rect 4331 10362 4337 10364
rect 4393 10362 4417 10364
rect 4473 10362 4497 10364
rect 4553 10362 4577 10364
rect 4633 10362 4639 10364
rect 4393 10310 4395 10362
rect 4575 10310 4577 10362
rect 4331 10308 4337 10310
rect 4393 10308 4417 10310
rect 4473 10308 4497 10310
rect 4553 10308 4577 10310
rect 4633 10308 4639 10310
rect 4331 10299 4639 10308
rect 5276 10266 5304 10610
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5276 10130 5304 10202
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4448 9518 4476 10066
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 5184 10010 5212 10066
rect 5460 10033 5488 10610
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5446 10024 5502 10033
rect 4540 9722 4568 9998
rect 4712 9988 4764 9994
rect 5184 9982 5446 10010
rect 5446 9959 5502 9968
rect 4712 9930 4764 9936
rect 4528 9716 4580 9722
rect 4528 9658 4580 9664
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4331 9276 4639 9285
rect 4331 9274 4337 9276
rect 4393 9274 4417 9276
rect 4473 9274 4497 9276
rect 4553 9274 4577 9276
rect 4633 9274 4639 9276
rect 4393 9222 4395 9274
rect 4575 9222 4577 9274
rect 4331 9220 4337 9222
rect 4393 9220 4417 9222
rect 4473 9220 4497 9222
rect 4553 9220 4577 9222
rect 4633 9220 4639 9222
rect 4331 9211 4639 9220
rect 4724 8634 4752 9930
rect 4991 9820 5299 9829
rect 4991 9818 4997 9820
rect 5053 9818 5077 9820
rect 5133 9818 5157 9820
rect 5213 9818 5237 9820
rect 5293 9818 5299 9820
rect 5053 9766 5055 9818
rect 5235 9766 5237 9818
rect 4991 9764 4997 9766
rect 5053 9764 5077 9766
rect 5133 9764 5157 9766
rect 5213 9764 5237 9766
rect 5293 9764 5299 9766
rect 4991 9755 5299 9764
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 5172 9376 5224 9382
rect 5224 9324 5396 9330
rect 5172 9318 5396 9324
rect 4816 9178 4844 9318
rect 5184 9302 5396 9318
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4991 8732 5299 8741
rect 4991 8730 4997 8732
rect 5053 8730 5077 8732
rect 5133 8730 5157 8732
rect 5213 8730 5237 8732
rect 5293 8730 5299 8732
rect 5053 8678 5055 8730
rect 5235 8678 5237 8730
rect 4991 8676 4997 8678
rect 5053 8676 5077 8678
rect 5133 8676 5157 8678
rect 5213 8676 5237 8678
rect 5293 8676 5299 8678
rect 4991 8667 5299 8676
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4712 8424 4764 8430
rect 4712 8366 4764 8372
rect 3436 8090 3464 8366
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3436 7546 3464 8026
rect 4172 7546 4200 8366
rect 4331 8188 4639 8197
rect 4331 8186 4337 8188
rect 4393 8186 4417 8188
rect 4473 8186 4497 8188
rect 4553 8186 4577 8188
rect 4633 8186 4639 8188
rect 4393 8134 4395 8186
rect 4575 8134 4577 8186
rect 4331 8132 4337 8134
rect 4393 8132 4417 8134
rect 4473 8132 4497 8134
rect 4553 8132 4577 8134
rect 4633 8132 4639 8134
rect 4331 8123 4639 8132
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4172 7041 4200 7346
rect 4158 7032 4214 7041
rect 4158 6967 4160 6976
rect 4212 6967 4214 6976
rect 4160 6938 4212 6944
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3896 5302 3924 5510
rect 2872 5296 2924 5302
rect 2872 5238 2924 5244
rect 3240 5296 3292 5302
rect 3240 5238 3292 5244
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 2077 4924 2385 4933
rect 2077 4922 2083 4924
rect 2139 4922 2163 4924
rect 2219 4922 2243 4924
rect 2299 4922 2323 4924
rect 2379 4922 2385 4924
rect 2139 4870 2141 4922
rect 2321 4870 2323 4922
rect 2077 4868 2083 4870
rect 2139 4868 2163 4870
rect 2219 4868 2243 4870
rect 2299 4868 2323 4870
rect 2379 4868 2385 4870
rect 2077 4859 2385 4868
rect 2884 4826 2912 5238
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2077 3836 2385 3845
rect 2077 3834 2083 3836
rect 2139 3834 2163 3836
rect 2219 3834 2243 3836
rect 2299 3834 2323 3836
rect 2379 3834 2385 3836
rect 2139 3782 2141 3834
rect 2321 3782 2323 3834
rect 2077 3780 2083 3782
rect 2139 3780 2163 3782
rect 2219 3780 2243 3782
rect 2299 3780 2323 3782
rect 2379 3780 2385 3782
rect 2077 3771 2385 3780
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 940 2848 992 2854
rect 938 2816 940 2825
rect 992 2816 994 2825
rect 938 2751 994 2760
rect 1504 2650 1532 2994
rect 2077 2748 2385 2757
rect 2077 2746 2083 2748
rect 2139 2746 2163 2748
rect 2219 2746 2243 2748
rect 2299 2746 2323 2748
rect 2379 2746 2385 2748
rect 2139 2694 2141 2746
rect 2321 2694 2323 2746
rect 2077 2692 2083 2694
rect 2139 2692 2163 2694
rect 2219 2692 2243 2694
rect 2299 2692 2323 2694
rect 2379 2692 2385 2694
rect 2077 2683 2385 2692
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 2424 2378 2452 4762
rect 2737 4380 3045 4389
rect 2737 4378 2743 4380
rect 2799 4378 2823 4380
rect 2879 4378 2903 4380
rect 2959 4378 2983 4380
rect 3039 4378 3045 4380
rect 2799 4326 2801 4378
rect 2981 4326 2983 4378
rect 2737 4324 2743 4326
rect 2799 4324 2823 4326
rect 2879 4324 2903 4326
rect 2959 4324 2983 4326
rect 3039 4324 3045 4326
rect 2737 4315 3045 4324
rect 2594 3496 2650 3505
rect 2594 3431 2650 3440
rect 2412 2372 2464 2378
rect 2412 2314 2464 2320
rect 20 2304 72 2310
rect 20 2246 72 2252
rect 32 800 60 2246
rect 2608 800 2636 3431
rect 2737 3292 3045 3301
rect 2737 3290 2743 3292
rect 2799 3290 2823 3292
rect 2879 3290 2903 3292
rect 2959 3290 2983 3292
rect 3039 3290 3045 3292
rect 2799 3238 2801 3290
rect 2981 3238 2983 3290
rect 2737 3236 2743 3238
rect 2799 3236 2823 3238
rect 2879 3236 2903 3238
rect 2959 3236 2983 3238
rect 3039 3236 3045 3238
rect 2737 3227 3045 3236
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2884 2514 2912 2790
rect 3344 2650 3372 5102
rect 3620 2922 3648 5102
rect 3698 4040 3754 4049
rect 3698 3975 3754 3984
rect 3712 3126 3740 3975
rect 4172 3505 4200 6666
rect 4264 6458 4292 7754
rect 4331 7100 4639 7109
rect 4331 7098 4337 7100
rect 4393 7098 4417 7100
rect 4473 7098 4497 7100
rect 4553 7098 4577 7100
rect 4633 7098 4639 7100
rect 4393 7046 4395 7098
rect 4575 7046 4577 7098
rect 4331 7044 4337 7046
rect 4393 7044 4417 7046
rect 4473 7044 4497 7046
rect 4553 7044 4577 7046
rect 4633 7044 4639 7046
rect 4331 7035 4639 7044
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4252 6316 4304 6322
rect 4252 6258 4304 6264
rect 4264 5642 4292 6258
rect 4331 6012 4639 6021
rect 4331 6010 4337 6012
rect 4393 6010 4417 6012
rect 4473 6010 4497 6012
rect 4553 6010 4577 6012
rect 4633 6010 4639 6012
rect 4393 5958 4395 6010
rect 4575 5958 4577 6010
rect 4331 5956 4337 5958
rect 4393 5956 4417 5958
rect 4473 5956 4497 5958
rect 4553 5956 4577 5958
rect 4633 5956 4639 5958
rect 4331 5947 4639 5956
rect 4724 5914 4752 8366
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7954 5212 8230
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7546 4936 7686
rect 4991 7644 5299 7653
rect 4991 7642 4997 7644
rect 5053 7642 5077 7644
rect 5133 7642 5157 7644
rect 5213 7642 5237 7644
rect 5293 7642 5299 7644
rect 5053 7590 5055 7642
rect 5235 7590 5237 7642
rect 4991 7588 4997 7590
rect 5053 7588 5077 7590
rect 5133 7588 5157 7590
rect 5213 7588 5237 7590
rect 5293 7588 5299 7590
rect 4991 7579 5299 7588
rect 5368 7546 5396 9302
rect 5460 7818 5488 9959
rect 5552 9382 5580 10406
rect 5644 9926 5672 10406
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 9722 5672 9862
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5828 9654 5856 10610
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5448 7812 5500 7818
rect 5448 7754 5500 7760
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 4816 6866 4844 7346
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4908 6798 4936 7142
rect 5552 7002 5580 7346
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6458 4936 6734
rect 4991 6556 5299 6565
rect 4991 6554 4997 6556
rect 5053 6554 5077 6556
rect 5133 6554 5157 6556
rect 5213 6554 5237 6556
rect 5293 6554 5299 6556
rect 5053 6502 5055 6554
rect 5235 6502 5237 6554
rect 4991 6500 4997 6502
rect 5053 6500 5077 6502
rect 5133 6500 5157 6502
rect 5213 6500 5237 6502
rect 5293 6500 5299 6502
rect 4991 6491 5299 6500
rect 5552 6458 5580 6938
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5092 6338 5120 6394
rect 4816 6322 5120 6338
rect 4804 6316 5120 6322
rect 4856 6310 5120 6316
rect 4804 6258 4856 6264
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4264 5370 4292 5578
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 4816 5166 4844 6258
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4908 5846 4936 6190
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 5092 5914 5120 6122
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 5736 5778 5764 7890
rect 5920 7886 5948 8230
rect 6288 7886 6316 8774
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6380 7818 6408 10406
rect 6585 10364 6893 10373
rect 6585 10362 6591 10364
rect 6647 10362 6671 10364
rect 6727 10362 6751 10364
rect 6807 10362 6831 10364
rect 6887 10362 6893 10364
rect 6647 10310 6649 10362
rect 6829 10310 6831 10362
rect 6585 10308 6591 10310
rect 6647 10308 6671 10310
rect 6727 10308 6751 10310
rect 6807 10308 6831 10310
rect 6887 10308 6893 10310
rect 6585 10299 6893 10308
rect 8839 10364 9147 10373
rect 8839 10362 8845 10364
rect 8901 10362 8925 10364
rect 8981 10362 9005 10364
rect 9061 10362 9085 10364
rect 9141 10362 9147 10364
rect 8901 10310 8903 10362
rect 9083 10310 9085 10362
rect 8839 10308 8845 10310
rect 8901 10308 8925 10310
rect 8981 10308 9005 10310
rect 9061 10308 9085 10310
rect 9141 10308 9147 10310
rect 8839 10299 9147 10308
rect 9324 10266 9352 10406
rect 9600 10266 9628 10406
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6472 8090 6500 10066
rect 8666 10024 8722 10033
rect 7104 9988 7156 9994
rect 8666 9959 8722 9968
rect 7104 9930 7156 9936
rect 6585 9276 6893 9285
rect 6585 9274 6591 9276
rect 6647 9274 6671 9276
rect 6727 9274 6751 9276
rect 6807 9274 6831 9276
rect 6887 9274 6893 9276
rect 6647 9222 6649 9274
rect 6829 9222 6831 9274
rect 6585 9220 6591 9222
rect 6647 9220 6671 9222
rect 6727 9220 6751 9222
rect 6807 9220 6831 9222
rect 6887 9220 6893 9222
rect 6585 9211 6893 9220
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6656 8362 6684 8910
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6585 8188 6893 8197
rect 6585 8186 6591 8188
rect 6647 8186 6671 8188
rect 6727 8186 6751 8188
rect 6807 8186 6831 8188
rect 6887 8186 6893 8188
rect 6647 8134 6649 8186
rect 6829 8134 6831 8186
rect 6585 8132 6591 8134
rect 6647 8132 6671 8134
rect 6727 8132 6751 8134
rect 6807 8132 6831 8134
rect 6887 8132 6893 8134
rect 6585 8123 6893 8132
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 6585 7100 6893 7109
rect 6585 7098 6591 7100
rect 6647 7098 6671 7100
rect 6727 7098 6751 7100
rect 6807 7098 6831 7100
rect 6887 7098 6893 7100
rect 6647 7046 6649 7098
rect 6829 7046 6831 7098
rect 6585 7044 6591 7046
rect 6647 7044 6671 7046
rect 6727 7044 6751 7046
rect 6807 7044 6831 7046
rect 6887 7044 6893 7046
rect 6585 7035 6893 7044
rect 6585 6012 6893 6021
rect 6585 6010 6591 6012
rect 6647 6010 6671 6012
rect 6727 6010 6751 6012
rect 6807 6010 6831 6012
rect 6887 6010 6893 6012
rect 6647 5958 6649 6010
rect 6829 5958 6831 6010
rect 6585 5956 6591 5958
rect 6647 5956 6671 5958
rect 6727 5956 6751 5958
rect 6807 5956 6831 5958
rect 6887 5956 6893 5958
rect 6585 5947 6893 5956
rect 6932 5794 6960 9114
rect 7116 8634 7144 9930
rect 8680 9926 8708 9959
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 7245 9820 7553 9829
rect 7245 9818 7251 9820
rect 7307 9818 7331 9820
rect 7387 9818 7411 9820
rect 7467 9818 7491 9820
rect 7547 9818 7553 9820
rect 7307 9766 7309 9818
rect 7489 9766 7491 9818
rect 7245 9764 7251 9766
rect 7307 9764 7331 9766
rect 7387 9764 7411 9766
rect 7467 9764 7491 9766
rect 7547 9764 7553 9766
rect 7245 9755 7553 9764
rect 7245 8732 7553 8741
rect 7245 8730 7251 8732
rect 7307 8730 7331 8732
rect 7387 8730 7411 8732
rect 7467 8730 7491 8732
rect 7547 8730 7553 8732
rect 7307 8678 7309 8730
rect 7489 8678 7491 8730
rect 7245 8676 7251 8678
rect 7307 8676 7331 8678
rect 7387 8676 7411 8678
rect 7467 8676 7491 8678
rect 7547 8676 7553 8678
rect 7245 8667 7553 8676
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 8208 8628 8260 8634
rect 8208 8570 8260 8576
rect 7116 7818 7144 8570
rect 8220 7970 8248 8570
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8404 8090 8432 8366
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8220 7942 8432 7970
rect 7104 7812 7156 7818
rect 7104 7754 7156 7760
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 7245 7644 7553 7653
rect 7245 7642 7251 7644
rect 7307 7642 7331 7644
rect 7387 7642 7411 7644
rect 7467 7642 7491 7644
rect 7547 7642 7553 7644
rect 7307 7590 7309 7642
rect 7489 7590 7491 7642
rect 7245 7588 7251 7590
rect 7307 7588 7331 7590
rect 7387 7588 7411 7590
rect 7467 7588 7491 7590
rect 7547 7588 7553 7590
rect 7245 7579 7553 7588
rect 8312 7410 8340 7686
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 7245 6556 7553 6565
rect 7245 6554 7251 6556
rect 7307 6554 7331 6556
rect 7387 6554 7411 6556
rect 7467 6554 7491 6556
rect 7547 6554 7553 6556
rect 7307 6502 7309 6554
rect 7489 6502 7491 6554
rect 7245 6500 7251 6502
rect 7307 6500 7331 6502
rect 7387 6500 7411 6502
rect 7467 6500 7491 6502
rect 7547 6500 7553 6502
rect 7245 6491 7553 6500
rect 8312 6474 8340 7346
rect 8220 6446 8340 6474
rect 8220 6390 8248 6446
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 5724 5772 5776 5778
rect 6932 5766 7144 5794
rect 5724 5714 5776 5720
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 4908 5302 4936 5510
rect 4991 5468 5299 5477
rect 4991 5466 4997 5468
rect 5053 5466 5077 5468
rect 5133 5466 5157 5468
rect 5213 5466 5237 5468
rect 5293 5466 5299 5468
rect 5053 5414 5055 5466
rect 5235 5414 5237 5466
rect 4991 5412 4997 5414
rect 5053 5412 5077 5414
rect 5133 5412 5157 5414
rect 5213 5412 5237 5414
rect 5293 5412 5299 5414
rect 4991 5403 5299 5412
rect 4896 5296 4948 5302
rect 4896 5238 4948 5244
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4331 4924 4639 4933
rect 4331 4922 4337 4924
rect 4393 4922 4417 4924
rect 4473 4922 4497 4924
rect 4553 4922 4577 4924
rect 4633 4922 4639 4924
rect 4393 4870 4395 4922
rect 4575 4870 4577 4922
rect 4331 4868 4337 4870
rect 4393 4868 4417 4870
rect 4473 4868 4497 4870
rect 4553 4868 4577 4870
rect 4633 4868 4639 4870
rect 4331 4859 4639 4868
rect 4331 3836 4639 3845
rect 4331 3834 4337 3836
rect 4393 3834 4417 3836
rect 4473 3834 4497 3836
rect 4553 3834 4577 3836
rect 4633 3834 4639 3836
rect 4393 3782 4395 3834
rect 4575 3782 4577 3834
rect 4331 3780 4337 3782
rect 4393 3780 4417 3782
rect 4473 3780 4497 3782
rect 4553 3780 4577 3782
rect 4633 3780 4639 3782
rect 4331 3771 4639 3780
rect 4158 3496 4214 3505
rect 4158 3431 4214 3440
rect 4908 3194 4936 5238
rect 4991 4380 5299 4389
rect 4991 4378 4997 4380
rect 5053 4378 5077 4380
rect 5133 4378 5157 4380
rect 5213 4378 5237 4380
rect 5293 4378 5299 4380
rect 5053 4326 5055 4378
rect 5235 4326 5237 4378
rect 4991 4324 4997 4326
rect 5053 4324 5077 4326
rect 5133 4324 5157 4326
rect 5213 4324 5237 4326
rect 5293 4324 5299 4326
rect 4991 4315 5299 4324
rect 4991 3292 5299 3301
rect 4991 3290 4997 3292
rect 5053 3290 5077 3292
rect 5133 3290 5157 3292
rect 5213 3290 5237 3292
rect 5293 3290 5299 3292
rect 5053 3238 5055 3290
rect 5235 3238 5237 3290
rect 4991 3236 4997 3238
rect 5053 3236 5077 3238
rect 5133 3236 5157 3238
rect 5213 3236 5237 3238
rect 5293 3236 5299 3238
rect 4991 3227 5299 3236
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5368 3126 5396 5510
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 4331 2748 4639 2757
rect 4331 2746 4337 2748
rect 4393 2746 4417 2748
rect 4473 2746 4497 2748
rect 4553 2746 4577 2748
rect 4633 2746 4639 2748
rect 4393 2694 4395 2746
rect 4575 2694 4577 2746
rect 4331 2692 4337 2694
rect 4393 2692 4417 2694
rect 4473 2692 4497 2694
rect 4553 2692 4577 2694
rect 4633 2692 4639 2694
rect 4331 2683 4639 2692
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 4724 2446 4752 2926
rect 6472 2650 6500 4966
rect 6585 4924 6893 4933
rect 6585 4922 6591 4924
rect 6647 4922 6671 4924
rect 6727 4922 6751 4924
rect 6807 4922 6831 4924
rect 6887 4922 6893 4924
rect 6647 4870 6649 4922
rect 6829 4870 6831 4922
rect 6585 4868 6591 4870
rect 6647 4868 6671 4870
rect 6727 4868 6751 4870
rect 6807 4868 6831 4870
rect 6887 4868 6893 4870
rect 6585 4859 6893 4868
rect 6585 3836 6893 3845
rect 6585 3834 6591 3836
rect 6647 3834 6671 3836
rect 6727 3834 6751 3836
rect 6807 3834 6831 3836
rect 6887 3834 6893 3836
rect 6647 3782 6649 3834
rect 6829 3782 6831 3834
rect 6585 3780 6591 3782
rect 6647 3780 6671 3782
rect 6727 3780 6751 3782
rect 6807 3780 6831 3782
rect 6887 3780 6893 3782
rect 6585 3771 6893 3780
rect 6932 3618 6960 5646
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7024 5370 7052 5510
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7116 5166 7144 5766
rect 7245 5468 7553 5477
rect 7245 5466 7251 5468
rect 7307 5466 7331 5468
rect 7387 5466 7411 5468
rect 7467 5466 7491 5468
rect 7547 5466 7553 5468
rect 7307 5414 7309 5466
rect 7489 5414 7491 5466
rect 7245 5412 7251 5414
rect 7307 5412 7331 5414
rect 7387 5412 7411 5414
rect 7467 5412 7491 5414
rect 7547 5412 7553 5414
rect 7245 5403 7553 5412
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 7116 4622 7144 5102
rect 7208 4826 7236 5170
rect 7300 5030 7328 5170
rect 7668 5166 7696 6054
rect 7852 5522 7880 6258
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 7760 5494 7880 5522
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7245 4380 7553 4389
rect 7245 4378 7251 4380
rect 7307 4378 7331 4380
rect 7387 4378 7411 4380
rect 7467 4378 7491 4380
rect 7547 4378 7553 4380
rect 7307 4326 7309 4378
rect 7489 4326 7491 4378
rect 7245 4324 7251 4326
rect 7307 4324 7331 4326
rect 7387 4324 7411 4326
rect 7467 4324 7491 4326
rect 7547 4324 7553 4326
rect 7245 4315 7553 4324
rect 6840 3590 6960 3618
rect 7668 3602 7696 4966
rect 7760 4622 7788 5494
rect 7944 5234 7972 6122
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 8220 5370 8248 6054
rect 8312 5914 8340 6122
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8404 5710 8432 7942
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7852 4826 7880 5170
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7656 3596 7708 3602
rect 6840 3534 6868 3590
rect 7656 3538 7708 3544
rect 8404 3534 8432 5646
rect 8588 5234 8616 5714
rect 8680 5710 8708 9862
rect 9499 9820 9807 9829
rect 9499 9818 9505 9820
rect 9561 9818 9585 9820
rect 9641 9818 9665 9820
rect 9721 9818 9745 9820
rect 9801 9818 9807 9820
rect 9561 9766 9563 9818
rect 9743 9766 9745 9818
rect 9499 9764 9505 9766
rect 9561 9764 9585 9766
rect 9641 9764 9665 9766
rect 9721 9764 9745 9766
rect 9801 9764 9807 9766
rect 9499 9755 9807 9764
rect 8839 9276 9147 9285
rect 8839 9274 8845 9276
rect 8901 9274 8925 9276
rect 8981 9274 9005 9276
rect 9061 9274 9085 9276
rect 9141 9274 9147 9276
rect 8901 9222 8903 9274
rect 9083 9222 9085 9274
rect 8839 9220 8845 9222
rect 8901 9220 8925 9222
rect 8981 9220 9005 9222
rect 9061 9220 9085 9222
rect 9141 9220 9147 9222
rect 8839 9211 9147 9220
rect 10140 8968 10192 8974
rect 10138 8936 10140 8945
rect 10192 8936 10194 8945
rect 10138 8871 10194 8880
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 8634 8892 8774
rect 9499 8732 9807 8741
rect 9499 8730 9505 8732
rect 9561 8730 9585 8732
rect 9641 8730 9665 8732
rect 9721 8730 9745 8732
rect 9801 8730 9807 8732
rect 9561 8678 9563 8730
rect 9743 8678 9745 8730
rect 9499 8676 9505 8678
rect 9561 8676 9585 8678
rect 9641 8676 9665 8678
rect 9721 8676 9745 8678
rect 9801 8676 9807 8678
rect 9499 8667 9807 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8839 8188 9147 8197
rect 8839 8186 8845 8188
rect 8901 8186 8925 8188
rect 8981 8186 9005 8188
rect 9061 8186 9085 8188
rect 9141 8186 9147 8188
rect 8901 8134 8903 8186
rect 9083 8134 9085 8186
rect 8839 8132 8845 8134
rect 8901 8132 8925 8134
rect 8981 8132 9005 8134
rect 9061 8132 9085 8134
rect 9141 8132 9147 8134
rect 8839 8123 9147 8132
rect 9499 7644 9807 7653
rect 9499 7642 9505 7644
rect 9561 7642 9585 7644
rect 9641 7642 9665 7644
rect 9721 7642 9745 7644
rect 9801 7642 9807 7644
rect 9561 7590 9563 7642
rect 9743 7590 9745 7642
rect 9499 7588 9505 7590
rect 9561 7588 9585 7590
rect 9641 7588 9665 7590
rect 9721 7588 9745 7590
rect 9801 7588 9807 7590
rect 9499 7579 9807 7588
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8772 6390 8800 7142
rect 8839 7100 9147 7109
rect 8839 7098 8845 7100
rect 8901 7098 8925 7100
rect 8981 7098 9005 7100
rect 9061 7098 9085 7100
rect 9141 7098 9147 7100
rect 8901 7046 8903 7098
rect 9083 7046 9085 7098
rect 8839 7044 8845 7046
rect 8901 7044 8925 7046
rect 8981 7044 9005 7046
rect 9061 7044 9085 7046
rect 9141 7044 9147 7046
rect 8839 7035 9147 7044
rect 9499 6556 9807 6565
rect 9499 6554 9505 6556
rect 9561 6554 9585 6556
rect 9641 6554 9665 6556
rect 9721 6554 9745 6556
rect 9801 6554 9807 6556
rect 9561 6502 9563 6554
rect 9743 6502 9745 6554
rect 9499 6500 9505 6502
rect 9561 6500 9585 6502
rect 9641 6500 9665 6502
rect 9721 6500 9745 6502
rect 9801 6500 9807 6502
rect 9499 6491 9807 6500
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8839 6012 9147 6021
rect 8839 6010 8845 6012
rect 8901 6010 8925 6012
rect 8981 6010 9005 6012
rect 9061 6010 9085 6012
rect 9141 6010 9147 6012
rect 8901 5958 8903 6010
rect 9083 5958 9085 6010
rect 8839 5956 8845 5958
rect 8901 5956 8925 5958
rect 8981 5956 9005 5958
rect 9061 5956 9085 5958
rect 9141 5956 9147 5958
rect 8839 5947 9147 5956
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8680 5302 8708 5646
rect 10048 5568 10100 5574
rect 10046 5536 10048 5545
rect 10100 5536 10102 5545
rect 9499 5468 9807 5477
rect 10046 5471 10102 5480
rect 9499 5466 9505 5468
rect 9561 5466 9585 5468
rect 9641 5466 9665 5468
rect 9721 5466 9745 5468
rect 9801 5466 9807 5468
rect 9561 5414 9563 5466
rect 9743 5414 9745 5466
rect 9499 5412 9505 5414
rect 9561 5412 9585 5414
rect 9641 5412 9665 5414
rect 9721 5412 9745 5414
rect 9801 5412 9807 5414
rect 9499 5403 9807 5412
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 6840 2990 6868 3470
rect 7245 3292 7553 3301
rect 7245 3290 7251 3292
rect 7307 3290 7331 3292
rect 7387 3290 7411 3292
rect 7467 3290 7491 3292
rect 7547 3290 7553 3292
rect 7307 3238 7309 3290
rect 7489 3238 7491 3290
rect 7245 3236 7251 3238
rect 7307 3236 7331 3238
rect 7387 3236 7411 3238
rect 7467 3236 7491 3238
rect 7547 3236 7553 3238
rect 7245 3227 7553 3236
rect 8404 3126 8432 3470
rect 8588 3194 8616 5170
rect 8668 5092 8720 5098
rect 8668 5034 8720 5040
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 6585 2748 6893 2757
rect 6585 2746 6591 2748
rect 6647 2746 6671 2748
rect 6727 2746 6751 2748
rect 6807 2746 6831 2748
rect 6887 2746 6893 2748
rect 6647 2694 6649 2746
rect 6829 2694 6831 2746
rect 6585 2692 6591 2694
rect 6647 2692 6671 2694
rect 6727 2692 6751 2694
rect 6807 2692 6831 2694
rect 6887 2692 6893 2694
rect 6585 2683 6893 2692
rect 8496 2650 8524 2926
rect 8680 2650 8708 5034
rect 8839 4924 9147 4933
rect 8839 4922 8845 4924
rect 8901 4922 8925 4924
rect 8981 4922 9005 4924
rect 9061 4922 9085 4924
rect 9141 4922 9147 4924
rect 8901 4870 8903 4922
rect 9083 4870 9085 4922
rect 8839 4868 8845 4870
rect 8901 4868 8925 4870
rect 8981 4868 9005 4870
rect 9061 4868 9085 4870
rect 9141 4868 9147 4870
rect 8839 4859 9147 4868
rect 9499 4380 9807 4389
rect 9499 4378 9505 4380
rect 9561 4378 9585 4380
rect 9641 4378 9665 4380
rect 9721 4378 9745 4380
rect 9801 4378 9807 4380
rect 9561 4326 9563 4378
rect 9743 4326 9745 4378
rect 9499 4324 9505 4326
rect 9561 4324 9585 4326
rect 9641 4324 9665 4326
rect 9721 4324 9745 4326
rect 9801 4324 9807 4326
rect 9499 4315 9807 4324
rect 8839 3836 9147 3845
rect 8839 3834 8845 3836
rect 8901 3834 8925 3836
rect 8981 3834 9005 3836
rect 9061 3834 9085 3836
rect 9141 3834 9147 3836
rect 8901 3782 8903 3834
rect 9083 3782 9085 3834
rect 8839 3780 8845 3782
rect 8901 3780 8925 3782
rect 8981 3780 9005 3782
rect 9061 3780 9085 3782
rect 9141 3780 9147 3782
rect 8839 3771 9147 3780
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 8772 3194 8800 3334
rect 9499 3292 9807 3301
rect 9499 3290 9505 3292
rect 9561 3290 9585 3292
rect 9641 3290 9665 3292
rect 9721 3290 9745 3292
rect 9801 3290 9807 3292
rect 9561 3238 9563 3290
rect 9743 3238 9745 3290
rect 9499 3236 9505 3238
rect 9561 3236 9585 3238
rect 9641 3236 9665 3238
rect 9721 3236 9745 3238
rect 9801 3236 9807 3238
rect 9499 3227 9807 3236
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 9680 2848 9732 2854
rect 9678 2816 9680 2825
rect 9732 2816 9734 2825
rect 8839 2748 9147 2757
rect 9678 2751 9734 2760
rect 8839 2746 8845 2748
rect 8901 2746 8925 2748
rect 8981 2746 9005 2748
rect 9061 2746 9085 2748
rect 9141 2746 9147 2748
rect 8901 2694 8903 2746
rect 9083 2694 9085 2746
rect 8839 2692 8845 2694
rect 8901 2692 8925 2694
rect 8981 2692 9005 2694
rect 9061 2692 9085 2694
rect 9141 2692 9147 2694
rect 8839 2683 9147 2692
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 2737 2204 3045 2213
rect 2737 2202 2743 2204
rect 2799 2202 2823 2204
rect 2879 2202 2903 2204
rect 2959 2202 2983 2204
rect 3039 2202 3045 2204
rect 2799 2150 2801 2202
rect 2981 2150 2983 2202
rect 2737 2148 2743 2150
rect 2799 2148 2823 2150
rect 2879 2148 2903 2150
rect 2959 2148 2983 2150
rect 3039 2148 3045 2150
rect 2737 2139 3045 2148
rect 4991 2204 5299 2213
rect 4991 2202 4997 2204
rect 5053 2202 5077 2204
rect 5133 2202 5157 2204
rect 5213 2202 5237 2204
rect 5293 2202 5299 2204
rect 5053 2150 5055 2202
rect 5235 2150 5237 2202
rect 4991 2148 4997 2150
rect 5053 2148 5077 2150
rect 5133 2148 5157 2150
rect 5213 2148 5237 2150
rect 5293 2148 5299 2150
rect 4991 2139 5299 2148
rect 5368 1170 5396 2246
rect 7245 2204 7553 2213
rect 7245 2202 7251 2204
rect 7307 2202 7331 2204
rect 7387 2202 7411 2204
rect 7467 2202 7491 2204
rect 7547 2202 7553 2204
rect 7307 2150 7309 2202
rect 7489 2150 7491 2202
rect 7245 2148 7251 2150
rect 7307 2148 7331 2150
rect 7387 2148 7411 2150
rect 7467 2148 7491 2150
rect 7547 2148 7553 2150
rect 7245 2139 7553 2148
rect 5184 1142 5396 1170
rect 5184 800 5212 1142
rect 8404 800 8432 2382
rect 9499 2204 9807 2213
rect 9499 2202 9505 2204
rect 9561 2202 9585 2204
rect 9641 2202 9665 2204
rect 9721 2202 9745 2204
rect 9801 2202 9807 2204
rect 9561 2150 9563 2202
rect 9743 2150 9745 2202
rect 9499 2148 9505 2150
rect 9561 2148 9585 2150
rect 9641 2148 9665 2150
rect 9721 2148 9745 2150
rect 9801 2148 9807 2150
rect 9499 2139 9807 2148
rect 10980 800 11008 2382
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 8390 0 8446 800
rect 10966 0 11022 800
<< via2 >>
rect 1950 11600 2006 11656
rect 2743 10906 2799 10908
rect 2823 10906 2879 10908
rect 2903 10906 2959 10908
rect 2983 10906 3039 10908
rect 2743 10854 2789 10906
rect 2789 10854 2799 10906
rect 2823 10854 2853 10906
rect 2853 10854 2865 10906
rect 2865 10854 2879 10906
rect 2903 10854 2917 10906
rect 2917 10854 2929 10906
rect 2929 10854 2959 10906
rect 2983 10854 2993 10906
rect 2993 10854 3039 10906
rect 2743 10852 2799 10854
rect 2823 10852 2879 10854
rect 2903 10852 2959 10854
rect 2983 10852 3039 10854
rect 4997 10906 5053 10908
rect 5077 10906 5133 10908
rect 5157 10906 5213 10908
rect 5237 10906 5293 10908
rect 4997 10854 5043 10906
rect 5043 10854 5053 10906
rect 5077 10854 5107 10906
rect 5107 10854 5119 10906
rect 5119 10854 5133 10906
rect 5157 10854 5171 10906
rect 5171 10854 5183 10906
rect 5183 10854 5213 10906
rect 5237 10854 5247 10906
rect 5247 10854 5293 10906
rect 4997 10852 5053 10854
rect 5077 10852 5133 10854
rect 5157 10852 5213 10854
rect 5237 10852 5293 10854
rect 9310 11600 9366 11656
rect 7251 10906 7307 10908
rect 7331 10906 7387 10908
rect 7411 10906 7467 10908
rect 7491 10906 7547 10908
rect 7251 10854 7297 10906
rect 7297 10854 7307 10906
rect 7331 10854 7361 10906
rect 7361 10854 7373 10906
rect 7373 10854 7387 10906
rect 7411 10854 7425 10906
rect 7425 10854 7437 10906
rect 7437 10854 7467 10906
rect 7491 10854 7501 10906
rect 7501 10854 7547 10906
rect 7251 10852 7307 10854
rect 7331 10852 7387 10854
rect 7411 10852 7467 10854
rect 7491 10852 7547 10854
rect 9505 10906 9561 10908
rect 9585 10906 9641 10908
rect 9665 10906 9721 10908
rect 9745 10906 9801 10908
rect 9505 10854 9551 10906
rect 9551 10854 9561 10906
rect 9585 10854 9615 10906
rect 9615 10854 9627 10906
rect 9627 10854 9641 10906
rect 9665 10854 9679 10906
rect 9679 10854 9691 10906
rect 9691 10854 9721 10906
rect 9745 10854 9755 10906
rect 9755 10854 9801 10906
rect 9505 10852 9561 10854
rect 9585 10852 9641 10854
rect 9665 10852 9721 10854
rect 9745 10852 9801 10854
rect 2083 10362 2139 10364
rect 2163 10362 2219 10364
rect 2243 10362 2299 10364
rect 2323 10362 2379 10364
rect 2083 10310 2129 10362
rect 2129 10310 2139 10362
rect 2163 10310 2193 10362
rect 2193 10310 2205 10362
rect 2205 10310 2219 10362
rect 2243 10310 2257 10362
rect 2257 10310 2269 10362
rect 2269 10310 2299 10362
rect 2323 10310 2333 10362
rect 2333 10310 2379 10362
rect 2083 10308 2139 10310
rect 2163 10308 2219 10310
rect 2243 10308 2299 10310
rect 2323 10308 2379 10310
rect 2743 9818 2799 9820
rect 2823 9818 2879 9820
rect 2903 9818 2959 9820
rect 2983 9818 3039 9820
rect 2743 9766 2789 9818
rect 2789 9766 2799 9818
rect 2823 9766 2853 9818
rect 2853 9766 2865 9818
rect 2865 9766 2879 9818
rect 2903 9766 2917 9818
rect 2917 9766 2929 9818
rect 2929 9766 2959 9818
rect 2983 9766 2993 9818
rect 2993 9766 3039 9818
rect 2743 9764 2799 9766
rect 2823 9764 2879 9766
rect 2903 9764 2959 9766
rect 2983 9764 3039 9766
rect 2083 9274 2139 9276
rect 2163 9274 2219 9276
rect 2243 9274 2299 9276
rect 2323 9274 2379 9276
rect 2083 9222 2129 9274
rect 2129 9222 2139 9274
rect 2163 9222 2193 9274
rect 2193 9222 2205 9274
rect 2205 9222 2219 9274
rect 2243 9222 2257 9274
rect 2257 9222 2269 9274
rect 2269 9222 2299 9274
rect 2323 9222 2333 9274
rect 2333 9222 2379 9274
rect 2083 9220 2139 9222
rect 2163 9220 2219 9222
rect 2243 9220 2299 9222
rect 2323 9220 2379 9222
rect 938 8880 994 8936
rect 2743 8730 2799 8732
rect 2823 8730 2879 8732
rect 2903 8730 2959 8732
rect 2983 8730 3039 8732
rect 2743 8678 2789 8730
rect 2789 8678 2799 8730
rect 2823 8678 2853 8730
rect 2853 8678 2865 8730
rect 2865 8678 2879 8730
rect 2903 8678 2917 8730
rect 2917 8678 2929 8730
rect 2929 8678 2959 8730
rect 2983 8678 2993 8730
rect 2993 8678 3039 8730
rect 2743 8676 2799 8678
rect 2823 8676 2879 8678
rect 2903 8676 2959 8678
rect 2983 8676 3039 8678
rect 2083 8186 2139 8188
rect 2163 8186 2219 8188
rect 2243 8186 2299 8188
rect 2323 8186 2379 8188
rect 2083 8134 2129 8186
rect 2129 8134 2139 8186
rect 2163 8134 2193 8186
rect 2193 8134 2205 8186
rect 2205 8134 2219 8186
rect 2243 8134 2257 8186
rect 2257 8134 2269 8186
rect 2269 8134 2299 8186
rect 2323 8134 2333 8186
rect 2333 8134 2379 8186
rect 2083 8132 2139 8134
rect 2163 8132 2219 8134
rect 2243 8132 2299 8134
rect 2323 8132 2379 8134
rect 2743 7642 2799 7644
rect 2823 7642 2879 7644
rect 2903 7642 2959 7644
rect 2983 7642 3039 7644
rect 2743 7590 2789 7642
rect 2789 7590 2799 7642
rect 2823 7590 2853 7642
rect 2853 7590 2865 7642
rect 2865 7590 2879 7642
rect 2903 7590 2917 7642
rect 2917 7590 2929 7642
rect 2929 7590 2959 7642
rect 2983 7590 2993 7642
rect 2993 7590 3039 7642
rect 2743 7588 2799 7590
rect 2823 7588 2879 7590
rect 2903 7588 2959 7590
rect 2983 7588 3039 7590
rect 2083 7098 2139 7100
rect 2163 7098 2219 7100
rect 2243 7098 2299 7100
rect 2323 7098 2379 7100
rect 2083 7046 2129 7098
rect 2129 7046 2139 7098
rect 2163 7046 2193 7098
rect 2193 7046 2205 7098
rect 2205 7046 2219 7098
rect 2243 7046 2257 7098
rect 2257 7046 2269 7098
rect 2269 7046 2299 7098
rect 2323 7046 2333 7098
rect 2333 7046 2379 7098
rect 2083 7044 2139 7046
rect 2163 7044 2219 7046
rect 2243 7044 2299 7046
rect 2323 7044 2379 7046
rect 2743 6554 2799 6556
rect 2823 6554 2879 6556
rect 2903 6554 2959 6556
rect 2983 6554 3039 6556
rect 2743 6502 2789 6554
rect 2789 6502 2799 6554
rect 2823 6502 2853 6554
rect 2853 6502 2865 6554
rect 2865 6502 2879 6554
rect 2903 6502 2917 6554
rect 2917 6502 2929 6554
rect 2929 6502 2959 6554
rect 2983 6502 2993 6554
rect 2993 6502 3039 6554
rect 2743 6500 2799 6502
rect 2823 6500 2879 6502
rect 2903 6500 2959 6502
rect 2983 6500 3039 6502
rect 2083 6010 2139 6012
rect 2163 6010 2219 6012
rect 2243 6010 2299 6012
rect 2323 6010 2379 6012
rect 2083 5958 2129 6010
rect 2129 5958 2139 6010
rect 2163 5958 2193 6010
rect 2193 5958 2205 6010
rect 2205 5958 2219 6010
rect 2243 5958 2257 6010
rect 2257 5958 2269 6010
rect 2269 5958 2299 6010
rect 2323 5958 2333 6010
rect 2333 5958 2379 6010
rect 2083 5956 2139 5958
rect 2163 5956 2219 5958
rect 2243 5956 2299 5958
rect 2323 5956 2379 5958
rect 1398 5480 1454 5536
rect 2743 5466 2799 5468
rect 2823 5466 2879 5468
rect 2903 5466 2959 5468
rect 2983 5466 3039 5468
rect 2743 5414 2789 5466
rect 2789 5414 2799 5466
rect 2823 5414 2853 5466
rect 2853 5414 2865 5466
rect 2865 5414 2879 5466
rect 2903 5414 2917 5466
rect 2917 5414 2929 5466
rect 2929 5414 2959 5466
rect 2983 5414 2993 5466
rect 2993 5414 3039 5466
rect 2743 5412 2799 5414
rect 2823 5412 2879 5414
rect 2903 5412 2959 5414
rect 2983 5412 3039 5414
rect 4337 10362 4393 10364
rect 4417 10362 4473 10364
rect 4497 10362 4553 10364
rect 4577 10362 4633 10364
rect 4337 10310 4383 10362
rect 4383 10310 4393 10362
rect 4417 10310 4447 10362
rect 4447 10310 4459 10362
rect 4459 10310 4473 10362
rect 4497 10310 4511 10362
rect 4511 10310 4523 10362
rect 4523 10310 4553 10362
rect 4577 10310 4587 10362
rect 4587 10310 4633 10362
rect 4337 10308 4393 10310
rect 4417 10308 4473 10310
rect 4497 10308 4553 10310
rect 4577 10308 4633 10310
rect 5446 9968 5502 10024
rect 4337 9274 4393 9276
rect 4417 9274 4473 9276
rect 4497 9274 4553 9276
rect 4577 9274 4633 9276
rect 4337 9222 4383 9274
rect 4383 9222 4393 9274
rect 4417 9222 4447 9274
rect 4447 9222 4459 9274
rect 4459 9222 4473 9274
rect 4497 9222 4511 9274
rect 4511 9222 4523 9274
rect 4523 9222 4553 9274
rect 4577 9222 4587 9274
rect 4587 9222 4633 9274
rect 4337 9220 4393 9222
rect 4417 9220 4473 9222
rect 4497 9220 4553 9222
rect 4577 9220 4633 9222
rect 4997 9818 5053 9820
rect 5077 9818 5133 9820
rect 5157 9818 5213 9820
rect 5237 9818 5293 9820
rect 4997 9766 5043 9818
rect 5043 9766 5053 9818
rect 5077 9766 5107 9818
rect 5107 9766 5119 9818
rect 5119 9766 5133 9818
rect 5157 9766 5171 9818
rect 5171 9766 5183 9818
rect 5183 9766 5213 9818
rect 5237 9766 5247 9818
rect 5247 9766 5293 9818
rect 4997 9764 5053 9766
rect 5077 9764 5133 9766
rect 5157 9764 5213 9766
rect 5237 9764 5293 9766
rect 4997 8730 5053 8732
rect 5077 8730 5133 8732
rect 5157 8730 5213 8732
rect 5237 8730 5293 8732
rect 4997 8678 5043 8730
rect 5043 8678 5053 8730
rect 5077 8678 5107 8730
rect 5107 8678 5119 8730
rect 5119 8678 5133 8730
rect 5157 8678 5171 8730
rect 5171 8678 5183 8730
rect 5183 8678 5213 8730
rect 5237 8678 5247 8730
rect 5247 8678 5293 8730
rect 4997 8676 5053 8678
rect 5077 8676 5133 8678
rect 5157 8676 5213 8678
rect 5237 8676 5293 8678
rect 4337 8186 4393 8188
rect 4417 8186 4473 8188
rect 4497 8186 4553 8188
rect 4577 8186 4633 8188
rect 4337 8134 4383 8186
rect 4383 8134 4393 8186
rect 4417 8134 4447 8186
rect 4447 8134 4459 8186
rect 4459 8134 4473 8186
rect 4497 8134 4511 8186
rect 4511 8134 4523 8186
rect 4523 8134 4553 8186
rect 4577 8134 4587 8186
rect 4587 8134 4633 8186
rect 4337 8132 4393 8134
rect 4417 8132 4473 8134
rect 4497 8132 4553 8134
rect 4577 8132 4633 8134
rect 4158 6996 4214 7032
rect 4158 6976 4160 6996
rect 4160 6976 4212 6996
rect 4212 6976 4214 6996
rect 2083 4922 2139 4924
rect 2163 4922 2219 4924
rect 2243 4922 2299 4924
rect 2323 4922 2379 4924
rect 2083 4870 2129 4922
rect 2129 4870 2139 4922
rect 2163 4870 2193 4922
rect 2193 4870 2205 4922
rect 2205 4870 2219 4922
rect 2243 4870 2257 4922
rect 2257 4870 2269 4922
rect 2269 4870 2299 4922
rect 2323 4870 2333 4922
rect 2333 4870 2379 4922
rect 2083 4868 2139 4870
rect 2163 4868 2219 4870
rect 2243 4868 2299 4870
rect 2323 4868 2379 4870
rect 2083 3834 2139 3836
rect 2163 3834 2219 3836
rect 2243 3834 2299 3836
rect 2323 3834 2379 3836
rect 2083 3782 2129 3834
rect 2129 3782 2139 3834
rect 2163 3782 2193 3834
rect 2193 3782 2205 3834
rect 2205 3782 2219 3834
rect 2243 3782 2257 3834
rect 2257 3782 2269 3834
rect 2269 3782 2299 3834
rect 2323 3782 2333 3834
rect 2333 3782 2379 3834
rect 2083 3780 2139 3782
rect 2163 3780 2219 3782
rect 2243 3780 2299 3782
rect 2323 3780 2379 3782
rect 938 2796 940 2816
rect 940 2796 992 2816
rect 992 2796 994 2816
rect 938 2760 994 2796
rect 2083 2746 2139 2748
rect 2163 2746 2219 2748
rect 2243 2746 2299 2748
rect 2323 2746 2379 2748
rect 2083 2694 2129 2746
rect 2129 2694 2139 2746
rect 2163 2694 2193 2746
rect 2193 2694 2205 2746
rect 2205 2694 2219 2746
rect 2243 2694 2257 2746
rect 2257 2694 2269 2746
rect 2269 2694 2299 2746
rect 2323 2694 2333 2746
rect 2333 2694 2379 2746
rect 2083 2692 2139 2694
rect 2163 2692 2219 2694
rect 2243 2692 2299 2694
rect 2323 2692 2379 2694
rect 2743 4378 2799 4380
rect 2823 4378 2879 4380
rect 2903 4378 2959 4380
rect 2983 4378 3039 4380
rect 2743 4326 2789 4378
rect 2789 4326 2799 4378
rect 2823 4326 2853 4378
rect 2853 4326 2865 4378
rect 2865 4326 2879 4378
rect 2903 4326 2917 4378
rect 2917 4326 2929 4378
rect 2929 4326 2959 4378
rect 2983 4326 2993 4378
rect 2993 4326 3039 4378
rect 2743 4324 2799 4326
rect 2823 4324 2879 4326
rect 2903 4324 2959 4326
rect 2983 4324 3039 4326
rect 2594 3440 2650 3496
rect 2743 3290 2799 3292
rect 2823 3290 2879 3292
rect 2903 3290 2959 3292
rect 2983 3290 3039 3292
rect 2743 3238 2789 3290
rect 2789 3238 2799 3290
rect 2823 3238 2853 3290
rect 2853 3238 2865 3290
rect 2865 3238 2879 3290
rect 2903 3238 2917 3290
rect 2917 3238 2929 3290
rect 2929 3238 2959 3290
rect 2983 3238 2993 3290
rect 2993 3238 3039 3290
rect 2743 3236 2799 3238
rect 2823 3236 2879 3238
rect 2903 3236 2959 3238
rect 2983 3236 3039 3238
rect 3698 3984 3754 4040
rect 4337 7098 4393 7100
rect 4417 7098 4473 7100
rect 4497 7098 4553 7100
rect 4577 7098 4633 7100
rect 4337 7046 4383 7098
rect 4383 7046 4393 7098
rect 4417 7046 4447 7098
rect 4447 7046 4459 7098
rect 4459 7046 4473 7098
rect 4497 7046 4511 7098
rect 4511 7046 4523 7098
rect 4523 7046 4553 7098
rect 4577 7046 4587 7098
rect 4587 7046 4633 7098
rect 4337 7044 4393 7046
rect 4417 7044 4473 7046
rect 4497 7044 4553 7046
rect 4577 7044 4633 7046
rect 4337 6010 4393 6012
rect 4417 6010 4473 6012
rect 4497 6010 4553 6012
rect 4577 6010 4633 6012
rect 4337 5958 4383 6010
rect 4383 5958 4393 6010
rect 4417 5958 4447 6010
rect 4447 5958 4459 6010
rect 4459 5958 4473 6010
rect 4497 5958 4511 6010
rect 4511 5958 4523 6010
rect 4523 5958 4553 6010
rect 4577 5958 4587 6010
rect 4587 5958 4633 6010
rect 4337 5956 4393 5958
rect 4417 5956 4473 5958
rect 4497 5956 4553 5958
rect 4577 5956 4633 5958
rect 4997 7642 5053 7644
rect 5077 7642 5133 7644
rect 5157 7642 5213 7644
rect 5237 7642 5293 7644
rect 4997 7590 5043 7642
rect 5043 7590 5053 7642
rect 5077 7590 5107 7642
rect 5107 7590 5119 7642
rect 5119 7590 5133 7642
rect 5157 7590 5171 7642
rect 5171 7590 5183 7642
rect 5183 7590 5213 7642
rect 5237 7590 5247 7642
rect 5247 7590 5293 7642
rect 4997 7588 5053 7590
rect 5077 7588 5133 7590
rect 5157 7588 5213 7590
rect 5237 7588 5293 7590
rect 4997 6554 5053 6556
rect 5077 6554 5133 6556
rect 5157 6554 5213 6556
rect 5237 6554 5293 6556
rect 4997 6502 5043 6554
rect 5043 6502 5053 6554
rect 5077 6502 5107 6554
rect 5107 6502 5119 6554
rect 5119 6502 5133 6554
rect 5157 6502 5171 6554
rect 5171 6502 5183 6554
rect 5183 6502 5213 6554
rect 5237 6502 5247 6554
rect 5247 6502 5293 6554
rect 4997 6500 5053 6502
rect 5077 6500 5133 6502
rect 5157 6500 5213 6502
rect 5237 6500 5293 6502
rect 6591 10362 6647 10364
rect 6671 10362 6727 10364
rect 6751 10362 6807 10364
rect 6831 10362 6887 10364
rect 6591 10310 6637 10362
rect 6637 10310 6647 10362
rect 6671 10310 6701 10362
rect 6701 10310 6713 10362
rect 6713 10310 6727 10362
rect 6751 10310 6765 10362
rect 6765 10310 6777 10362
rect 6777 10310 6807 10362
rect 6831 10310 6841 10362
rect 6841 10310 6887 10362
rect 6591 10308 6647 10310
rect 6671 10308 6727 10310
rect 6751 10308 6807 10310
rect 6831 10308 6887 10310
rect 8845 10362 8901 10364
rect 8925 10362 8981 10364
rect 9005 10362 9061 10364
rect 9085 10362 9141 10364
rect 8845 10310 8891 10362
rect 8891 10310 8901 10362
rect 8925 10310 8955 10362
rect 8955 10310 8967 10362
rect 8967 10310 8981 10362
rect 9005 10310 9019 10362
rect 9019 10310 9031 10362
rect 9031 10310 9061 10362
rect 9085 10310 9095 10362
rect 9095 10310 9141 10362
rect 8845 10308 8901 10310
rect 8925 10308 8981 10310
rect 9005 10308 9061 10310
rect 9085 10308 9141 10310
rect 8666 9968 8722 10024
rect 6591 9274 6647 9276
rect 6671 9274 6727 9276
rect 6751 9274 6807 9276
rect 6831 9274 6887 9276
rect 6591 9222 6637 9274
rect 6637 9222 6647 9274
rect 6671 9222 6701 9274
rect 6701 9222 6713 9274
rect 6713 9222 6727 9274
rect 6751 9222 6765 9274
rect 6765 9222 6777 9274
rect 6777 9222 6807 9274
rect 6831 9222 6841 9274
rect 6841 9222 6887 9274
rect 6591 9220 6647 9222
rect 6671 9220 6727 9222
rect 6751 9220 6807 9222
rect 6831 9220 6887 9222
rect 6591 8186 6647 8188
rect 6671 8186 6727 8188
rect 6751 8186 6807 8188
rect 6831 8186 6887 8188
rect 6591 8134 6637 8186
rect 6637 8134 6647 8186
rect 6671 8134 6701 8186
rect 6701 8134 6713 8186
rect 6713 8134 6727 8186
rect 6751 8134 6765 8186
rect 6765 8134 6777 8186
rect 6777 8134 6807 8186
rect 6831 8134 6841 8186
rect 6841 8134 6887 8186
rect 6591 8132 6647 8134
rect 6671 8132 6727 8134
rect 6751 8132 6807 8134
rect 6831 8132 6887 8134
rect 6591 7098 6647 7100
rect 6671 7098 6727 7100
rect 6751 7098 6807 7100
rect 6831 7098 6887 7100
rect 6591 7046 6637 7098
rect 6637 7046 6647 7098
rect 6671 7046 6701 7098
rect 6701 7046 6713 7098
rect 6713 7046 6727 7098
rect 6751 7046 6765 7098
rect 6765 7046 6777 7098
rect 6777 7046 6807 7098
rect 6831 7046 6841 7098
rect 6841 7046 6887 7098
rect 6591 7044 6647 7046
rect 6671 7044 6727 7046
rect 6751 7044 6807 7046
rect 6831 7044 6887 7046
rect 6591 6010 6647 6012
rect 6671 6010 6727 6012
rect 6751 6010 6807 6012
rect 6831 6010 6887 6012
rect 6591 5958 6637 6010
rect 6637 5958 6647 6010
rect 6671 5958 6701 6010
rect 6701 5958 6713 6010
rect 6713 5958 6727 6010
rect 6751 5958 6765 6010
rect 6765 5958 6777 6010
rect 6777 5958 6807 6010
rect 6831 5958 6841 6010
rect 6841 5958 6887 6010
rect 6591 5956 6647 5958
rect 6671 5956 6727 5958
rect 6751 5956 6807 5958
rect 6831 5956 6887 5958
rect 7251 9818 7307 9820
rect 7331 9818 7387 9820
rect 7411 9818 7467 9820
rect 7491 9818 7547 9820
rect 7251 9766 7297 9818
rect 7297 9766 7307 9818
rect 7331 9766 7361 9818
rect 7361 9766 7373 9818
rect 7373 9766 7387 9818
rect 7411 9766 7425 9818
rect 7425 9766 7437 9818
rect 7437 9766 7467 9818
rect 7491 9766 7501 9818
rect 7501 9766 7547 9818
rect 7251 9764 7307 9766
rect 7331 9764 7387 9766
rect 7411 9764 7467 9766
rect 7491 9764 7547 9766
rect 7251 8730 7307 8732
rect 7331 8730 7387 8732
rect 7411 8730 7467 8732
rect 7491 8730 7547 8732
rect 7251 8678 7297 8730
rect 7297 8678 7307 8730
rect 7331 8678 7361 8730
rect 7361 8678 7373 8730
rect 7373 8678 7387 8730
rect 7411 8678 7425 8730
rect 7425 8678 7437 8730
rect 7437 8678 7467 8730
rect 7491 8678 7501 8730
rect 7501 8678 7547 8730
rect 7251 8676 7307 8678
rect 7331 8676 7387 8678
rect 7411 8676 7467 8678
rect 7491 8676 7547 8678
rect 7251 7642 7307 7644
rect 7331 7642 7387 7644
rect 7411 7642 7467 7644
rect 7491 7642 7547 7644
rect 7251 7590 7297 7642
rect 7297 7590 7307 7642
rect 7331 7590 7361 7642
rect 7361 7590 7373 7642
rect 7373 7590 7387 7642
rect 7411 7590 7425 7642
rect 7425 7590 7437 7642
rect 7437 7590 7467 7642
rect 7491 7590 7501 7642
rect 7501 7590 7547 7642
rect 7251 7588 7307 7590
rect 7331 7588 7387 7590
rect 7411 7588 7467 7590
rect 7491 7588 7547 7590
rect 7251 6554 7307 6556
rect 7331 6554 7387 6556
rect 7411 6554 7467 6556
rect 7491 6554 7547 6556
rect 7251 6502 7297 6554
rect 7297 6502 7307 6554
rect 7331 6502 7361 6554
rect 7361 6502 7373 6554
rect 7373 6502 7387 6554
rect 7411 6502 7425 6554
rect 7425 6502 7437 6554
rect 7437 6502 7467 6554
rect 7491 6502 7501 6554
rect 7501 6502 7547 6554
rect 7251 6500 7307 6502
rect 7331 6500 7387 6502
rect 7411 6500 7467 6502
rect 7491 6500 7547 6502
rect 4997 5466 5053 5468
rect 5077 5466 5133 5468
rect 5157 5466 5213 5468
rect 5237 5466 5293 5468
rect 4997 5414 5043 5466
rect 5043 5414 5053 5466
rect 5077 5414 5107 5466
rect 5107 5414 5119 5466
rect 5119 5414 5133 5466
rect 5157 5414 5171 5466
rect 5171 5414 5183 5466
rect 5183 5414 5213 5466
rect 5237 5414 5247 5466
rect 5247 5414 5293 5466
rect 4997 5412 5053 5414
rect 5077 5412 5133 5414
rect 5157 5412 5213 5414
rect 5237 5412 5293 5414
rect 4337 4922 4393 4924
rect 4417 4922 4473 4924
rect 4497 4922 4553 4924
rect 4577 4922 4633 4924
rect 4337 4870 4383 4922
rect 4383 4870 4393 4922
rect 4417 4870 4447 4922
rect 4447 4870 4459 4922
rect 4459 4870 4473 4922
rect 4497 4870 4511 4922
rect 4511 4870 4523 4922
rect 4523 4870 4553 4922
rect 4577 4870 4587 4922
rect 4587 4870 4633 4922
rect 4337 4868 4393 4870
rect 4417 4868 4473 4870
rect 4497 4868 4553 4870
rect 4577 4868 4633 4870
rect 4337 3834 4393 3836
rect 4417 3834 4473 3836
rect 4497 3834 4553 3836
rect 4577 3834 4633 3836
rect 4337 3782 4383 3834
rect 4383 3782 4393 3834
rect 4417 3782 4447 3834
rect 4447 3782 4459 3834
rect 4459 3782 4473 3834
rect 4497 3782 4511 3834
rect 4511 3782 4523 3834
rect 4523 3782 4553 3834
rect 4577 3782 4587 3834
rect 4587 3782 4633 3834
rect 4337 3780 4393 3782
rect 4417 3780 4473 3782
rect 4497 3780 4553 3782
rect 4577 3780 4633 3782
rect 4158 3440 4214 3496
rect 4997 4378 5053 4380
rect 5077 4378 5133 4380
rect 5157 4378 5213 4380
rect 5237 4378 5293 4380
rect 4997 4326 5043 4378
rect 5043 4326 5053 4378
rect 5077 4326 5107 4378
rect 5107 4326 5119 4378
rect 5119 4326 5133 4378
rect 5157 4326 5171 4378
rect 5171 4326 5183 4378
rect 5183 4326 5213 4378
rect 5237 4326 5247 4378
rect 5247 4326 5293 4378
rect 4997 4324 5053 4326
rect 5077 4324 5133 4326
rect 5157 4324 5213 4326
rect 5237 4324 5293 4326
rect 4997 3290 5053 3292
rect 5077 3290 5133 3292
rect 5157 3290 5213 3292
rect 5237 3290 5293 3292
rect 4997 3238 5043 3290
rect 5043 3238 5053 3290
rect 5077 3238 5107 3290
rect 5107 3238 5119 3290
rect 5119 3238 5133 3290
rect 5157 3238 5171 3290
rect 5171 3238 5183 3290
rect 5183 3238 5213 3290
rect 5237 3238 5247 3290
rect 5247 3238 5293 3290
rect 4997 3236 5053 3238
rect 5077 3236 5133 3238
rect 5157 3236 5213 3238
rect 5237 3236 5293 3238
rect 4337 2746 4393 2748
rect 4417 2746 4473 2748
rect 4497 2746 4553 2748
rect 4577 2746 4633 2748
rect 4337 2694 4383 2746
rect 4383 2694 4393 2746
rect 4417 2694 4447 2746
rect 4447 2694 4459 2746
rect 4459 2694 4473 2746
rect 4497 2694 4511 2746
rect 4511 2694 4523 2746
rect 4523 2694 4553 2746
rect 4577 2694 4587 2746
rect 4587 2694 4633 2746
rect 4337 2692 4393 2694
rect 4417 2692 4473 2694
rect 4497 2692 4553 2694
rect 4577 2692 4633 2694
rect 6591 4922 6647 4924
rect 6671 4922 6727 4924
rect 6751 4922 6807 4924
rect 6831 4922 6887 4924
rect 6591 4870 6637 4922
rect 6637 4870 6647 4922
rect 6671 4870 6701 4922
rect 6701 4870 6713 4922
rect 6713 4870 6727 4922
rect 6751 4870 6765 4922
rect 6765 4870 6777 4922
rect 6777 4870 6807 4922
rect 6831 4870 6841 4922
rect 6841 4870 6887 4922
rect 6591 4868 6647 4870
rect 6671 4868 6727 4870
rect 6751 4868 6807 4870
rect 6831 4868 6887 4870
rect 6591 3834 6647 3836
rect 6671 3834 6727 3836
rect 6751 3834 6807 3836
rect 6831 3834 6887 3836
rect 6591 3782 6637 3834
rect 6637 3782 6647 3834
rect 6671 3782 6701 3834
rect 6701 3782 6713 3834
rect 6713 3782 6727 3834
rect 6751 3782 6765 3834
rect 6765 3782 6777 3834
rect 6777 3782 6807 3834
rect 6831 3782 6841 3834
rect 6841 3782 6887 3834
rect 6591 3780 6647 3782
rect 6671 3780 6727 3782
rect 6751 3780 6807 3782
rect 6831 3780 6887 3782
rect 7251 5466 7307 5468
rect 7331 5466 7387 5468
rect 7411 5466 7467 5468
rect 7491 5466 7547 5468
rect 7251 5414 7297 5466
rect 7297 5414 7307 5466
rect 7331 5414 7361 5466
rect 7361 5414 7373 5466
rect 7373 5414 7387 5466
rect 7411 5414 7425 5466
rect 7425 5414 7437 5466
rect 7437 5414 7467 5466
rect 7491 5414 7501 5466
rect 7501 5414 7547 5466
rect 7251 5412 7307 5414
rect 7331 5412 7387 5414
rect 7411 5412 7467 5414
rect 7491 5412 7547 5414
rect 7251 4378 7307 4380
rect 7331 4378 7387 4380
rect 7411 4378 7467 4380
rect 7491 4378 7547 4380
rect 7251 4326 7297 4378
rect 7297 4326 7307 4378
rect 7331 4326 7361 4378
rect 7361 4326 7373 4378
rect 7373 4326 7387 4378
rect 7411 4326 7425 4378
rect 7425 4326 7437 4378
rect 7437 4326 7467 4378
rect 7491 4326 7501 4378
rect 7501 4326 7547 4378
rect 7251 4324 7307 4326
rect 7331 4324 7387 4326
rect 7411 4324 7467 4326
rect 7491 4324 7547 4326
rect 9505 9818 9561 9820
rect 9585 9818 9641 9820
rect 9665 9818 9721 9820
rect 9745 9818 9801 9820
rect 9505 9766 9551 9818
rect 9551 9766 9561 9818
rect 9585 9766 9615 9818
rect 9615 9766 9627 9818
rect 9627 9766 9641 9818
rect 9665 9766 9679 9818
rect 9679 9766 9691 9818
rect 9691 9766 9721 9818
rect 9745 9766 9755 9818
rect 9755 9766 9801 9818
rect 9505 9764 9561 9766
rect 9585 9764 9641 9766
rect 9665 9764 9721 9766
rect 9745 9764 9801 9766
rect 8845 9274 8901 9276
rect 8925 9274 8981 9276
rect 9005 9274 9061 9276
rect 9085 9274 9141 9276
rect 8845 9222 8891 9274
rect 8891 9222 8901 9274
rect 8925 9222 8955 9274
rect 8955 9222 8967 9274
rect 8967 9222 8981 9274
rect 9005 9222 9019 9274
rect 9019 9222 9031 9274
rect 9031 9222 9061 9274
rect 9085 9222 9095 9274
rect 9095 9222 9141 9274
rect 8845 9220 8901 9222
rect 8925 9220 8981 9222
rect 9005 9220 9061 9222
rect 9085 9220 9141 9222
rect 10138 8916 10140 8936
rect 10140 8916 10192 8936
rect 10192 8916 10194 8936
rect 10138 8880 10194 8916
rect 9505 8730 9561 8732
rect 9585 8730 9641 8732
rect 9665 8730 9721 8732
rect 9745 8730 9801 8732
rect 9505 8678 9551 8730
rect 9551 8678 9561 8730
rect 9585 8678 9615 8730
rect 9615 8678 9627 8730
rect 9627 8678 9641 8730
rect 9665 8678 9679 8730
rect 9679 8678 9691 8730
rect 9691 8678 9721 8730
rect 9745 8678 9755 8730
rect 9755 8678 9801 8730
rect 9505 8676 9561 8678
rect 9585 8676 9641 8678
rect 9665 8676 9721 8678
rect 9745 8676 9801 8678
rect 8845 8186 8901 8188
rect 8925 8186 8981 8188
rect 9005 8186 9061 8188
rect 9085 8186 9141 8188
rect 8845 8134 8891 8186
rect 8891 8134 8901 8186
rect 8925 8134 8955 8186
rect 8955 8134 8967 8186
rect 8967 8134 8981 8186
rect 9005 8134 9019 8186
rect 9019 8134 9031 8186
rect 9031 8134 9061 8186
rect 9085 8134 9095 8186
rect 9095 8134 9141 8186
rect 8845 8132 8901 8134
rect 8925 8132 8981 8134
rect 9005 8132 9061 8134
rect 9085 8132 9141 8134
rect 9505 7642 9561 7644
rect 9585 7642 9641 7644
rect 9665 7642 9721 7644
rect 9745 7642 9801 7644
rect 9505 7590 9551 7642
rect 9551 7590 9561 7642
rect 9585 7590 9615 7642
rect 9615 7590 9627 7642
rect 9627 7590 9641 7642
rect 9665 7590 9679 7642
rect 9679 7590 9691 7642
rect 9691 7590 9721 7642
rect 9745 7590 9755 7642
rect 9755 7590 9801 7642
rect 9505 7588 9561 7590
rect 9585 7588 9641 7590
rect 9665 7588 9721 7590
rect 9745 7588 9801 7590
rect 8845 7098 8901 7100
rect 8925 7098 8981 7100
rect 9005 7098 9061 7100
rect 9085 7098 9141 7100
rect 8845 7046 8891 7098
rect 8891 7046 8901 7098
rect 8925 7046 8955 7098
rect 8955 7046 8967 7098
rect 8967 7046 8981 7098
rect 9005 7046 9019 7098
rect 9019 7046 9031 7098
rect 9031 7046 9061 7098
rect 9085 7046 9095 7098
rect 9095 7046 9141 7098
rect 8845 7044 8901 7046
rect 8925 7044 8981 7046
rect 9005 7044 9061 7046
rect 9085 7044 9141 7046
rect 9505 6554 9561 6556
rect 9585 6554 9641 6556
rect 9665 6554 9721 6556
rect 9745 6554 9801 6556
rect 9505 6502 9551 6554
rect 9551 6502 9561 6554
rect 9585 6502 9615 6554
rect 9615 6502 9627 6554
rect 9627 6502 9641 6554
rect 9665 6502 9679 6554
rect 9679 6502 9691 6554
rect 9691 6502 9721 6554
rect 9745 6502 9755 6554
rect 9755 6502 9801 6554
rect 9505 6500 9561 6502
rect 9585 6500 9641 6502
rect 9665 6500 9721 6502
rect 9745 6500 9801 6502
rect 8845 6010 8901 6012
rect 8925 6010 8981 6012
rect 9005 6010 9061 6012
rect 9085 6010 9141 6012
rect 8845 5958 8891 6010
rect 8891 5958 8901 6010
rect 8925 5958 8955 6010
rect 8955 5958 8967 6010
rect 8967 5958 8981 6010
rect 9005 5958 9019 6010
rect 9019 5958 9031 6010
rect 9031 5958 9061 6010
rect 9085 5958 9095 6010
rect 9095 5958 9141 6010
rect 8845 5956 8901 5958
rect 8925 5956 8981 5958
rect 9005 5956 9061 5958
rect 9085 5956 9141 5958
rect 10046 5516 10048 5536
rect 10048 5516 10100 5536
rect 10100 5516 10102 5536
rect 10046 5480 10102 5516
rect 9505 5466 9561 5468
rect 9585 5466 9641 5468
rect 9665 5466 9721 5468
rect 9745 5466 9801 5468
rect 9505 5414 9551 5466
rect 9551 5414 9561 5466
rect 9585 5414 9615 5466
rect 9615 5414 9627 5466
rect 9627 5414 9641 5466
rect 9665 5414 9679 5466
rect 9679 5414 9691 5466
rect 9691 5414 9721 5466
rect 9745 5414 9755 5466
rect 9755 5414 9801 5466
rect 9505 5412 9561 5414
rect 9585 5412 9641 5414
rect 9665 5412 9721 5414
rect 9745 5412 9801 5414
rect 7251 3290 7307 3292
rect 7331 3290 7387 3292
rect 7411 3290 7467 3292
rect 7491 3290 7547 3292
rect 7251 3238 7297 3290
rect 7297 3238 7307 3290
rect 7331 3238 7361 3290
rect 7361 3238 7373 3290
rect 7373 3238 7387 3290
rect 7411 3238 7425 3290
rect 7425 3238 7437 3290
rect 7437 3238 7467 3290
rect 7491 3238 7501 3290
rect 7501 3238 7547 3290
rect 7251 3236 7307 3238
rect 7331 3236 7387 3238
rect 7411 3236 7467 3238
rect 7491 3236 7547 3238
rect 6591 2746 6647 2748
rect 6671 2746 6727 2748
rect 6751 2746 6807 2748
rect 6831 2746 6887 2748
rect 6591 2694 6637 2746
rect 6637 2694 6647 2746
rect 6671 2694 6701 2746
rect 6701 2694 6713 2746
rect 6713 2694 6727 2746
rect 6751 2694 6765 2746
rect 6765 2694 6777 2746
rect 6777 2694 6807 2746
rect 6831 2694 6841 2746
rect 6841 2694 6887 2746
rect 6591 2692 6647 2694
rect 6671 2692 6727 2694
rect 6751 2692 6807 2694
rect 6831 2692 6887 2694
rect 8845 4922 8901 4924
rect 8925 4922 8981 4924
rect 9005 4922 9061 4924
rect 9085 4922 9141 4924
rect 8845 4870 8891 4922
rect 8891 4870 8901 4922
rect 8925 4870 8955 4922
rect 8955 4870 8967 4922
rect 8967 4870 8981 4922
rect 9005 4870 9019 4922
rect 9019 4870 9031 4922
rect 9031 4870 9061 4922
rect 9085 4870 9095 4922
rect 9095 4870 9141 4922
rect 8845 4868 8901 4870
rect 8925 4868 8981 4870
rect 9005 4868 9061 4870
rect 9085 4868 9141 4870
rect 9505 4378 9561 4380
rect 9585 4378 9641 4380
rect 9665 4378 9721 4380
rect 9745 4378 9801 4380
rect 9505 4326 9551 4378
rect 9551 4326 9561 4378
rect 9585 4326 9615 4378
rect 9615 4326 9627 4378
rect 9627 4326 9641 4378
rect 9665 4326 9679 4378
rect 9679 4326 9691 4378
rect 9691 4326 9721 4378
rect 9745 4326 9755 4378
rect 9755 4326 9801 4378
rect 9505 4324 9561 4326
rect 9585 4324 9641 4326
rect 9665 4324 9721 4326
rect 9745 4324 9801 4326
rect 8845 3834 8901 3836
rect 8925 3834 8981 3836
rect 9005 3834 9061 3836
rect 9085 3834 9141 3836
rect 8845 3782 8891 3834
rect 8891 3782 8901 3834
rect 8925 3782 8955 3834
rect 8955 3782 8967 3834
rect 8967 3782 8981 3834
rect 9005 3782 9019 3834
rect 9019 3782 9031 3834
rect 9031 3782 9061 3834
rect 9085 3782 9095 3834
rect 9095 3782 9141 3834
rect 8845 3780 8901 3782
rect 8925 3780 8981 3782
rect 9005 3780 9061 3782
rect 9085 3780 9141 3782
rect 9505 3290 9561 3292
rect 9585 3290 9641 3292
rect 9665 3290 9721 3292
rect 9745 3290 9801 3292
rect 9505 3238 9551 3290
rect 9551 3238 9561 3290
rect 9585 3238 9615 3290
rect 9615 3238 9627 3290
rect 9627 3238 9641 3290
rect 9665 3238 9679 3290
rect 9679 3238 9691 3290
rect 9691 3238 9721 3290
rect 9745 3238 9755 3290
rect 9755 3238 9801 3290
rect 9505 3236 9561 3238
rect 9585 3236 9641 3238
rect 9665 3236 9721 3238
rect 9745 3236 9801 3238
rect 9678 2796 9680 2816
rect 9680 2796 9732 2816
rect 9732 2796 9734 2816
rect 9678 2760 9734 2796
rect 8845 2746 8901 2748
rect 8925 2746 8981 2748
rect 9005 2746 9061 2748
rect 9085 2746 9141 2748
rect 8845 2694 8891 2746
rect 8891 2694 8901 2746
rect 8925 2694 8955 2746
rect 8955 2694 8967 2746
rect 8967 2694 8981 2746
rect 9005 2694 9019 2746
rect 9019 2694 9031 2746
rect 9031 2694 9061 2746
rect 9085 2694 9095 2746
rect 9095 2694 9141 2746
rect 8845 2692 8901 2694
rect 8925 2692 8981 2694
rect 9005 2692 9061 2694
rect 9085 2692 9141 2694
rect 2743 2202 2799 2204
rect 2823 2202 2879 2204
rect 2903 2202 2959 2204
rect 2983 2202 3039 2204
rect 2743 2150 2789 2202
rect 2789 2150 2799 2202
rect 2823 2150 2853 2202
rect 2853 2150 2865 2202
rect 2865 2150 2879 2202
rect 2903 2150 2917 2202
rect 2917 2150 2929 2202
rect 2929 2150 2959 2202
rect 2983 2150 2993 2202
rect 2993 2150 3039 2202
rect 2743 2148 2799 2150
rect 2823 2148 2879 2150
rect 2903 2148 2959 2150
rect 2983 2148 3039 2150
rect 4997 2202 5053 2204
rect 5077 2202 5133 2204
rect 5157 2202 5213 2204
rect 5237 2202 5293 2204
rect 4997 2150 5043 2202
rect 5043 2150 5053 2202
rect 5077 2150 5107 2202
rect 5107 2150 5119 2202
rect 5119 2150 5133 2202
rect 5157 2150 5171 2202
rect 5171 2150 5183 2202
rect 5183 2150 5213 2202
rect 5237 2150 5247 2202
rect 5247 2150 5293 2202
rect 4997 2148 5053 2150
rect 5077 2148 5133 2150
rect 5157 2148 5213 2150
rect 5237 2148 5293 2150
rect 7251 2202 7307 2204
rect 7331 2202 7387 2204
rect 7411 2202 7467 2204
rect 7491 2202 7547 2204
rect 7251 2150 7297 2202
rect 7297 2150 7307 2202
rect 7331 2150 7361 2202
rect 7361 2150 7373 2202
rect 7373 2150 7387 2202
rect 7411 2150 7425 2202
rect 7425 2150 7437 2202
rect 7437 2150 7467 2202
rect 7491 2150 7501 2202
rect 7501 2150 7547 2202
rect 7251 2148 7307 2150
rect 7331 2148 7387 2150
rect 7411 2148 7467 2150
rect 7491 2148 7547 2150
rect 9505 2202 9561 2204
rect 9585 2202 9641 2204
rect 9665 2202 9721 2204
rect 9745 2202 9801 2204
rect 9505 2150 9551 2202
rect 9551 2150 9561 2202
rect 9585 2150 9615 2202
rect 9615 2150 9627 2202
rect 9627 2150 9641 2202
rect 9665 2150 9679 2202
rect 9679 2150 9691 2202
rect 9691 2150 9721 2202
rect 9745 2150 9755 2202
rect 9755 2150 9801 2202
rect 9505 2148 9561 2150
rect 9585 2148 9641 2150
rect 9665 2148 9721 2150
rect 9745 2148 9801 2150
<< metal3 >>
rect 0 11658 800 11688
rect 1945 11658 2011 11661
rect 0 11656 2011 11658
rect 0 11600 1950 11656
rect 2006 11600 2011 11656
rect 0 11598 2011 11600
rect 0 11568 800 11598
rect 1945 11595 2011 11598
rect 9305 11658 9371 11661
rect 10495 11658 11295 11688
rect 9305 11656 11295 11658
rect 9305 11600 9310 11656
rect 9366 11600 11295 11656
rect 9305 11598 11295 11600
rect 9305 11595 9371 11598
rect 10495 11568 11295 11598
rect 2733 10912 3049 10913
rect 2733 10848 2739 10912
rect 2803 10848 2819 10912
rect 2883 10848 2899 10912
rect 2963 10848 2979 10912
rect 3043 10848 3049 10912
rect 2733 10847 3049 10848
rect 4987 10912 5303 10913
rect 4987 10848 4993 10912
rect 5057 10848 5073 10912
rect 5137 10848 5153 10912
rect 5217 10848 5233 10912
rect 5297 10848 5303 10912
rect 4987 10847 5303 10848
rect 7241 10912 7557 10913
rect 7241 10848 7247 10912
rect 7311 10848 7327 10912
rect 7391 10848 7407 10912
rect 7471 10848 7487 10912
rect 7551 10848 7557 10912
rect 7241 10847 7557 10848
rect 9495 10912 9811 10913
rect 9495 10848 9501 10912
rect 9565 10848 9581 10912
rect 9645 10848 9661 10912
rect 9725 10848 9741 10912
rect 9805 10848 9811 10912
rect 9495 10847 9811 10848
rect 2073 10368 2389 10369
rect 2073 10304 2079 10368
rect 2143 10304 2159 10368
rect 2223 10304 2239 10368
rect 2303 10304 2319 10368
rect 2383 10304 2389 10368
rect 2073 10303 2389 10304
rect 4327 10368 4643 10369
rect 4327 10304 4333 10368
rect 4397 10304 4413 10368
rect 4477 10304 4493 10368
rect 4557 10304 4573 10368
rect 4637 10304 4643 10368
rect 4327 10303 4643 10304
rect 6581 10368 6897 10369
rect 6581 10304 6587 10368
rect 6651 10304 6667 10368
rect 6731 10304 6747 10368
rect 6811 10304 6827 10368
rect 6891 10304 6897 10368
rect 6581 10303 6897 10304
rect 8835 10368 9151 10369
rect 8835 10304 8841 10368
rect 8905 10304 8921 10368
rect 8985 10304 9001 10368
rect 9065 10304 9081 10368
rect 9145 10304 9151 10368
rect 8835 10303 9151 10304
rect 5441 10026 5507 10029
rect 8661 10026 8727 10029
rect 5441 10024 8727 10026
rect 5441 9968 5446 10024
rect 5502 9968 8666 10024
rect 8722 9968 8727 10024
rect 5441 9966 8727 9968
rect 5441 9963 5507 9966
rect 8661 9963 8727 9966
rect 2733 9824 3049 9825
rect 2733 9760 2739 9824
rect 2803 9760 2819 9824
rect 2883 9760 2899 9824
rect 2963 9760 2979 9824
rect 3043 9760 3049 9824
rect 2733 9759 3049 9760
rect 4987 9824 5303 9825
rect 4987 9760 4993 9824
rect 5057 9760 5073 9824
rect 5137 9760 5153 9824
rect 5217 9760 5233 9824
rect 5297 9760 5303 9824
rect 4987 9759 5303 9760
rect 7241 9824 7557 9825
rect 7241 9760 7247 9824
rect 7311 9760 7327 9824
rect 7391 9760 7407 9824
rect 7471 9760 7487 9824
rect 7551 9760 7557 9824
rect 7241 9759 7557 9760
rect 9495 9824 9811 9825
rect 9495 9760 9501 9824
rect 9565 9760 9581 9824
rect 9645 9760 9661 9824
rect 9725 9760 9741 9824
rect 9805 9760 9811 9824
rect 9495 9759 9811 9760
rect 2073 9280 2389 9281
rect 2073 9216 2079 9280
rect 2143 9216 2159 9280
rect 2223 9216 2239 9280
rect 2303 9216 2319 9280
rect 2383 9216 2389 9280
rect 2073 9215 2389 9216
rect 4327 9280 4643 9281
rect 4327 9216 4333 9280
rect 4397 9216 4413 9280
rect 4477 9216 4493 9280
rect 4557 9216 4573 9280
rect 4637 9216 4643 9280
rect 4327 9215 4643 9216
rect 6581 9280 6897 9281
rect 6581 9216 6587 9280
rect 6651 9216 6667 9280
rect 6731 9216 6747 9280
rect 6811 9216 6827 9280
rect 6891 9216 6897 9280
rect 6581 9215 6897 9216
rect 8835 9280 9151 9281
rect 8835 9216 8841 9280
rect 8905 9216 8921 9280
rect 8985 9216 9001 9280
rect 9065 9216 9081 9280
rect 9145 9216 9151 9280
rect 8835 9215 9151 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 10133 8938 10199 8941
rect 10495 8938 11295 8968
rect 10133 8936 11295 8938
rect 10133 8880 10138 8936
rect 10194 8880 11295 8936
rect 10133 8878 11295 8880
rect 10133 8875 10199 8878
rect 10495 8848 11295 8878
rect 2733 8736 3049 8737
rect 2733 8672 2739 8736
rect 2803 8672 2819 8736
rect 2883 8672 2899 8736
rect 2963 8672 2979 8736
rect 3043 8672 3049 8736
rect 2733 8671 3049 8672
rect 4987 8736 5303 8737
rect 4987 8672 4993 8736
rect 5057 8672 5073 8736
rect 5137 8672 5153 8736
rect 5217 8672 5233 8736
rect 5297 8672 5303 8736
rect 4987 8671 5303 8672
rect 7241 8736 7557 8737
rect 7241 8672 7247 8736
rect 7311 8672 7327 8736
rect 7391 8672 7407 8736
rect 7471 8672 7487 8736
rect 7551 8672 7557 8736
rect 7241 8671 7557 8672
rect 9495 8736 9811 8737
rect 9495 8672 9501 8736
rect 9565 8672 9581 8736
rect 9645 8672 9661 8736
rect 9725 8672 9741 8736
rect 9805 8672 9811 8736
rect 9495 8671 9811 8672
rect 2073 8192 2389 8193
rect 2073 8128 2079 8192
rect 2143 8128 2159 8192
rect 2223 8128 2239 8192
rect 2303 8128 2319 8192
rect 2383 8128 2389 8192
rect 2073 8127 2389 8128
rect 4327 8192 4643 8193
rect 4327 8128 4333 8192
rect 4397 8128 4413 8192
rect 4477 8128 4493 8192
rect 4557 8128 4573 8192
rect 4637 8128 4643 8192
rect 4327 8127 4643 8128
rect 6581 8192 6897 8193
rect 6581 8128 6587 8192
rect 6651 8128 6667 8192
rect 6731 8128 6747 8192
rect 6811 8128 6827 8192
rect 6891 8128 6897 8192
rect 6581 8127 6897 8128
rect 8835 8192 9151 8193
rect 8835 8128 8841 8192
rect 8905 8128 8921 8192
rect 8985 8128 9001 8192
rect 9065 8128 9081 8192
rect 9145 8128 9151 8192
rect 8835 8127 9151 8128
rect 2733 7648 3049 7649
rect 2733 7584 2739 7648
rect 2803 7584 2819 7648
rect 2883 7584 2899 7648
rect 2963 7584 2979 7648
rect 3043 7584 3049 7648
rect 2733 7583 3049 7584
rect 4987 7648 5303 7649
rect 4987 7584 4993 7648
rect 5057 7584 5073 7648
rect 5137 7584 5153 7648
rect 5217 7584 5233 7648
rect 5297 7584 5303 7648
rect 4987 7583 5303 7584
rect 7241 7648 7557 7649
rect 7241 7584 7247 7648
rect 7311 7584 7327 7648
rect 7391 7584 7407 7648
rect 7471 7584 7487 7648
rect 7551 7584 7557 7648
rect 7241 7583 7557 7584
rect 9495 7648 9811 7649
rect 9495 7584 9501 7648
rect 9565 7584 9581 7648
rect 9645 7584 9661 7648
rect 9725 7584 9741 7648
rect 9805 7584 9811 7648
rect 9495 7583 9811 7584
rect 2073 7104 2389 7105
rect 2073 7040 2079 7104
rect 2143 7040 2159 7104
rect 2223 7040 2239 7104
rect 2303 7040 2319 7104
rect 2383 7040 2389 7104
rect 2073 7039 2389 7040
rect 4327 7104 4643 7105
rect 4327 7040 4333 7104
rect 4397 7040 4413 7104
rect 4477 7040 4493 7104
rect 4557 7040 4573 7104
rect 4637 7040 4643 7104
rect 4327 7039 4643 7040
rect 6581 7104 6897 7105
rect 6581 7040 6587 7104
rect 6651 7040 6667 7104
rect 6731 7040 6747 7104
rect 6811 7040 6827 7104
rect 6891 7040 6897 7104
rect 6581 7039 6897 7040
rect 8835 7104 9151 7105
rect 8835 7040 8841 7104
rect 8905 7040 8921 7104
rect 8985 7040 9001 7104
rect 9065 7040 9081 7104
rect 9145 7040 9151 7104
rect 8835 7039 9151 7040
rect 4153 7036 4219 7037
rect 4102 6972 4108 7036
rect 4172 7034 4219 7036
rect 4172 7032 4264 7034
rect 4214 6976 4264 7032
rect 4172 6974 4264 6976
rect 4172 6972 4219 6974
rect 4153 6971 4219 6972
rect 2733 6560 3049 6561
rect 2733 6496 2739 6560
rect 2803 6496 2819 6560
rect 2883 6496 2899 6560
rect 2963 6496 2979 6560
rect 3043 6496 3049 6560
rect 2733 6495 3049 6496
rect 4987 6560 5303 6561
rect 4987 6496 4993 6560
rect 5057 6496 5073 6560
rect 5137 6496 5153 6560
rect 5217 6496 5233 6560
rect 5297 6496 5303 6560
rect 4987 6495 5303 6496
rect 7241 6560 7557 6561
rect 7241 6496 7247 6560
rect 7311 6496 7327 6560
rect 7391 6496 7407 6560
rect 7471 6496 7487 6560
rect 7551 6496 7557 6560
rect 7241 6495 7557 6496
rect 9495 6560 9811 6561
rect 9495 6496 9501 6560
rect 9565 6496 9581 6560
rect 9645 6496 9661 6560
rect 9725 6496 9741 6560
rect 9805 6496 9811 6560
rect 9495 6495 9811 6496
rect 2073 6016 2389 6017
rect 2073 5952 2079 6016
rect 2143 5952 2159 6016
rect 2223 5952 2239 6016
rect 2303 5952 2319 6016
rect 2383 5952 2389 6016
rect 2073 5951 2389 5952
rect 4327 6016 4643 6017
rect 4327 5952 4333 6016
rect 4397 5952 4413 6016
rect 4477 5952 4493 6016
rect 4557 5952 4573 6016
rect 4637 5952 4643 6016
rect 4327 5951 4643 5952
rect 6581 6016 6897 6017
rect 6581 5952 6587 6016
rect 6651 5952 6667 6016
rect 6731 5952 6747 6016
rect 6811 5952 6827 6016
rect 6891 5952 6897 6016
rect 6581 5951 6897 5952
rect 8835 6016 9151 6017
rect 8835 5952 8841 6016
rect 8905 5952 8921 6016
rect 8985 5952 9001 6016
rect 9065 5952 9081 6016
rect 9145 5952 9151 6016
rect 8835 5951 9151 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 10041 5538 10107 5541
rect 10495 5538 11295 5568
rect 10041 5536 11295 5538
rect 10041 5480 10046 5536
rect 10102 5480 11295 5536
rect 10041 5478 11295 5480
rect 10041 5475 10107 5478
rect 2733 5472 3049 5473
rect 2733 5408 2739 5472
rect 2803 5408 2819 5472
rect 2883 5408 2899 5472
rect 2963 5408 2979 5472
rect 3043 5408 3049 5472
rect 2733 5407 3049 5408
rect 4987 5472 5303 5473
rect 4987 5408 4993 5472
rect 5057 5408 5073 5472
rect 5137 5408 5153 5472
rect 5217 5408 5233 5472
rect 5297 5408 5303 5472
rect 4987 5407 5303 5408
rect 7241 5472 7557 5473
rect 7241 5408 7247 5472
rect 7311 5408 7327 5472
rect 7391 5408 7407 5472
rect 7471 5408 7487 5472
rect 7551 5408 7557 5472
rect 7241 5407 7557 5408
rect 9495 5472 9811 5473
rect 9495 5408 9501 5472
rect 9565 5408 9581 5472
rect 9645 5408 9661 5472
rect 9725 5408 9741 5472
rect 9805 5408 9811 5472
rect 10495 5448 11295 5478
rect 9495 5407 9811 5408
rect 2073 4928 2389 4929
rect 2073 4864 2079 4928
rect 2143 4864 2159 4928
rect 2223 4864 2239 4928
rect 2303 4864 2319 4928
rect 2383 4864 2389 4928
rect 2073 4863 2389 4864
rect 4327 4928 4643 4929
rect 4327 4864 4333 4928
rect 4397 4864 4413 4928
rect 4477 4864 4493 4928
rect 4557 4864 4573 4928
rect 4637 4864 4643 4928
rect 4327 4863 4643 4864
rect 6581 4928 6897 4929
rect 6581 4864 6587 4928
rect 6651 4864 6667 4928
rect 6731 4864 6747 4928
rect 6811 4864 6827 4928
rect 6891 4864 6897 4928
rect 6581 4863 6897 4864
rect 8835 4928 9151 4929
rect 8835 4864 8841 4928
rect 8905 4864 8921 4928
rect 8985 4864 9001 4928
rect 9065 4864 9081 4928
rect 9145 4864 9151 4928
rect 8835 4863 9151 4864
rect 2733 4384 3049 4385
rect 2733 4320 2739 4384
rect 2803 4320 2819 4384
rect 2883 4320 2899 4384
rect 2963 4320 2979 4384
rect 3043 4320 3049 4384
rect 2733 4319 3049 4320
rect 4987 4384 5303 4385
rect 4987 4320 4993 4384
rect 5057 4320 5073 4384
rect 5137 4320 5153 4384
rect 5217 4320 5233 4384
rect 5297 4320 5303 4384
rect 4987 4319 5303 4320
rect 7241 4384 7557 4385
rect 7241 4320 7247 4384
rect 7311 4320 7327 4384
rect 7391 4320 7407 4384
rect 7471 4320 7487 4384
rect 7551 4320 7557 4384
rect 7241 4319 7557 4320
rect 9495 4384 9811 4385
rect 9495 4320 9501 4384
rect 9565 4320 9581 4384
rect 9645 4320 9661 4384
rect 9725 4320 9741 4384
rect 9805 4320 9811 4384
rect 9495 4319 9811 4320
rect 3693 4042 3759 4045
rect 4102 4042 4108 4044
rect 3693 4040 4108 4042
rect 3693 3984 3698 4040
rect 3754 3984 4108 4040
rect 3693 3982 4108 3984
rect 3693 3979 3759 3982
rect 4102 3980 4108 3982
rect 4172 3980 4178 4044
rect 2073 3840 2389 3841
rect 2073 3776 2079 3840
rect 2143 3776 2159 3840
rect 2223 3776 2239 3840
rect 2303 3776 2319 3840
rect 2383 3776 2389 3840
rect 2073 3775 2389 3776
rect 4327 3840 4643 3841
rect 4327 3776 4333 3840
rect 4397 3776 4413 3840
rect 4477 3776 4493 3840
rect 4557 3776 4573 3840
rect 4637 3776 4643 3840
rect 4327 3775 4643 3776
rect 6581 3840 6897 3841
rect 6581 3776 6587 3840
rect 6651 3776 6667 3840
rect 6731 3776 6747 3840
rect 6811 3776 6827 3840
rect 6891 3776 6897 3840
rect 6581 3775 6897 3776
rect 8835 3840 9151 3841
rect 8835 3776 8841 3840
rect 8905 3776 8921 3840
rect 8985 3776 9001 3840
rect 9065 3776 9081 3840
rect 9145 3776 9151 3840
rect 8835 3775 9151 3776
rect 2589 3498 2655 3501
rect 4153 3498 4219 3501
rect 2589 3496 4219 3498
rect 2589 3440 2594 3496
rect 2650 3440 4158 3496
rect 4214 3440 4219 3496
rect 2589 3438 4219 3440
rect 2589 3435 2655 3438
rect 4153 3435 4219 3438
rect 2733 3296 3049 3297
rect 2733 3232 2739 3296
rect 2803 3232 2819 3296
rect 2883 3232 2899 3296
rect 2963 3232 2979 3296
rect 3043 3232 3049 3296
rect 2733 3231 3049 3232
rect 4987 3296 5303 3297
rect 4987 3232 4993 3296
rect 5057 3232 5073 3296
rect 5137 3232 5153 3296
rect 5217 3232 5233 3296
rect 5297 3232 5303 3296
rect 4987 3231 5303 3232
rect 7241 3296 7557 3297
rect 7241 3232 7247 3296
rect 7311 3232 7327 3296
rect 7391 3232 7407 3296
rect 7471 3232 7487 3296
rect 7551 3232 7557 3296
rect 7241 3231 7557 3232
rect 9495 3296 9811 3297
rect 9495 3232 9501 3296
rect 9565 3232 9581 3296
rect 9645 3232 9661 3296
rect 9725 3232 9741 3296
rect 9805 3232 9811 3296
rect 9495 3231 9811 3232
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 9673 2818 9739 2821
rect 10495 2818 11295 2848
rect 9673 2816 11295 2818
rect 9673 2760 9678 2816
rect 9734 2760 11295 2816
rect 9673 2758 11295 2760
rect 9673 2755 9739 2758
rect 2073 2752 2389 2753
rect 2073 2688 2079 2752
rect 2143 2688 2159 2752
rect 2223 2688 2239 2752
rect 2303 2688 2319 2752
rect 2383 2688 2389 2752
rect 2073 2687 2389 2688
rect 4327 2752 4643 2753
rect 4327 2688 4333 2752
rect 4397 2688 4413 2752
rect 4477 2688 4493 2752
rect 4557 2688 4573 2752
rect 4637 2688 4643 2752
rect 4327 2687 4643 2688
rect 6581 2752 6897 2753
rect 6581 2688 6587 2752
rect 6651 2688 6667 2752
rect 6731 2688 6747 2752
rect 6811 2688 6827 2752
rect 6891 2688 6897 2752
rect 6581 2687 6897 2688
rect 8835 2752 9151 2753
rect 8835 2688 8841 2752
rect 8905 2688 8921 2752
rect 8985 2688 9001 2752
rect 9065 2688 9081 2752
rect 9145 2688 9151 2752
rect 10495 2728 11295 2758
rect 8835 2687 9151 2688
rect 2733 2208 3049 2209
rect 2733 2144 2739 2208
rect 2803 2144 2819 2208
rect 2883 2144 2899 2208
rect 2963 2144 2979 2208
rect 3043 2144 3049 2208
rect 2733 2143 3049 2144
rect 4987 2208 5303 2209
rect 4987 2144 4993 2208
rect 5057 2144 5073 2208
rect 5137 2144 5153 2208
rect 5217 2144 5233 2208
rect 5297 2144 5303 2208
rect 4987 2143 5303 2144
rect 7241 2208 7557 2209
rect 7241 2144 7247 2208
rect 7311 2144 7327 2208
rect 7391 2144 7407 2208
rect 7471 2144 7487 2208
rect 7551 2144 7557 2208
rect 7241 2143 7557 2144
rect 9495 2208 9811 2209
rect 9495 2144 9501 2208
rect 9565 2144 9581 2208
rect 9645 2144 9661 2208
rect 9725 2144 9741 2208
rect 9805 2144 9811 2208
rect 9495 2143 9811 2144
<< via3 >>
rect 2739 10908 2803 10912
rect 2739 10852 2743 10908
rect 2743 10852 2799 10908
rect 2799 10852 2803 10908
rect 2739 10848 2803 10852
rect 2819 10908 2883 10912
rect 2819 10852 2823 10908
rect 2823 10852 2879 10908
rect 2879 10852 2883 10908
rect 2819 10848 2883 10852
rect 2899 10908 2963 10912
rect 2899 10852 2903 10908
rect 2903 10852 2959 10908
rect 2959 10852 2963 10908
rect 2899 10848 2963 10852
rect 2979 10908 3043 10912
rect 2979 10852 2983 10908
rect 2983 10852 3039 10908
rect 3039 10852 3043 10908
rect 2979 10848 3043 10852
rect 4993 10908 5057 10912
rect 4993 10852 4997 10908
rect 4997 10852 5053 10908
rect 5053 10852 5057 10908
rect 4993 10848 5057 10852
rect 5073 10908 5137 10912
rect 5073 10852 5077 10908
rect 5077 10852 5133 10908
rect 5133 10852 5137 10908
rect 5073 10848 5137 10852
rect 5153 10908 5217 10912
rect 5153 10852 5157 10908
rect 5157 10852 5213 10908
rect 5213 10852 5217 10908
rect 5153 10848 5217 10852
rect 5233 10908 5297 10912
rect 5233 10852 5237 10908
rect 5237 10852 5293 10908
rect 5293 10852 5297 10908
rect 5233 10848 5297 10852
rect 7247 10908 7311 10912
rect 7247 10852 7251 10908
rect 7251 10852 7307 10908
rect 7307 10852 7311 10908
rect 7247 10848 7311 10852
rect 7327 10908 7391 10912
rect 7327 10852 7331 10908
rect 7331 10852 7387 10908
rect 7387 10852 7391 10908
rect 7327 10848 7391 10852
rect 7407 10908 7471 10912
rect 7407 10852 7411 10908
rect 7411 10852 7467 10908
rect 7467 10852 7471 10908
rect 7407 10848 7471 10852
rect 7487 10908 7551 10912
rect 7487 10852 7491 10908
rect 7491 10852 7547 10908
rect 7547 10852 7551 10908
rect 7487 10848 7551 10852
rect 9501 10908 9565 10912
rect 9501 10852 9505 10908
rect 9505 10852 9561 10908
rect 9561 10852 9565 10908
rect 9501 10848 9565 10852
rect 9581 10908 9645 10912
rect 9581 10852 9585 10908
rect 9585 10852 9641 10908
rect 9641 10852 9645 10908
rect 9581 10848 9645 10852
rect 9661 10908 9725 10912
rect 9661 10852 9665 10908
rect 9665 10852 9721 10908
rect 9721 10852 9725 10908
rect 9661 10848 9725 10852
rect 9741 10908 9805 10912
rect 9741 10852 9745 10908
rect 9745 10852 9801 10908
rect 9801 10852 9805 10908
rect 9741 10848 9805 10852
rect 2079 10364 2143 10368
rect 2079 10308 2083 10364
rect 2083 10308 2139 10364
rect 2139 10308 2143 10364
rect 2079 10304 2143 10308
rect 2159 10364 2223 10368
rect 2159 10308 2163 10364
rect 2163 10308 2219 10364
rect 2219 10308 2223 10364
rect 2159 10304 2223 10308
rect 2239 10364 2303 10368
rect 2239 10308 2243 10364
rect 2243 10308 2299 10364
rect 2299 10308 2303 10364
rect 2239 10304 2303 10308
rect 2319 10364 2383 10368
rect 2319 10308 2323 10364
rect 2323 10308 2379 10364
rect 2379 10308 2383 10364
rect 2319 10304 2383 10308
rect 4333 10364 4397 10368
rect 4333 10308 4337 10364
rect 4337 10308 4393 10364
rect 4393 10308 4397 10364
rect 4333 10304 4397 10308
rect 4413 10364 4477 10368
rect 4413 10308 4417 10364
rect 4417 10308 4473 10364
rect 4473 10308 4477 10364
rect 4413 10304 4477 10308
rect 4493 10364 4557 10368
rect 4493 10308 4497 10364
rect 4497 10308 4553 10364
rect 4553 10308 4557 10364
rect 4493 10304 4557 10308
rect 4573 10364 4637 10368
rect 4573 10308 4577 10364
rect 4577 10308 4633 10364
rect 4633 10308 4637 10364
rect 4573 10304 4637 10308
rect 6587 10364 6651 10368
rect 6587 10308 6591 10364
rect 6591 10308 6647 10364
rect 6647 10308 6651 10364
rect 6587 10304 6651 10308
rect 6667 10364 6731 10368
rect 6667 10308 6671 10364
rect 6671 10308 6727 10364
rect 6727 10308 6731 10364
rect 6667 10304 6731 10308
rect 6747 10364 6811 10368
rect 6747 10308 6751 10364
rect 6751 10308 6807 10364
rect 6807 10308 6811 10364
rect 6747 10304 6811 10308
rect 6827 10364 6891 10368
rect 6827 10308 6831 10364
rect 6831 10308 6887 10364
rect 6887 10308 6891 10364
rect 6827 10304 6891 10308
rect 8841 10364 8905 10368
rect 8841 10308 8845 10364
rect 8845 10308 8901 10364
rect 8901 10308 8905 10364
rect 8841 10304 8905 10308
rect 8921 10364 8985 10368
rect 8921 10308 8925 10364
rect 8925 10308 8981 10364
rect 8981 10308 8985 10364
rect 8921 10304 8985 10308
rect 9001 10364 9065 10368
rect 9001 10308 9005 10364
rect 9005 10308 9061 10364
rect 9061 10308 9065 10364
rect 9001 10304 9065 10308
rect 9081 10364 9145 10368
rect 9081 10308 9085 10364
rect 9085 10308 9141 10364
rect 9141 10308 9145 10364
rect 9081 10304 9145 10308
rect 2739 9820 2803 9824
rect 2739 9764 2743 9820
rect 2743 9764 2799 9820
rect 2799 9764 2803 9820
rect 2739 9760 2803 9764
rect 2819 9820 2883 9824
rect 2819 9764 2823 9820
rect 2823 9764 2879 9820
rect 2879 9764 2883 9820
rect 2819 9760 2883 9764
rect 2899 9820 2963 9824
rect 2899 9764 2903 9820
rect 2903 9764 2959 9820
rect 2959 9764 2963 9820
rect 2899 9760 2963 9764
rect 2979 9820 3043 9824
rect 2979 9764 2983 9820
rect 2983 9764 3039 9820
rect 3039 9764 3043 9820
rect 2979 9760 3043 9764
rect 4993 9820 5057 9824
rect 4993 9764 4997 9820
rect 4997 9764 5053 9820
rect 5053 9764 5057 9820
rect 4993 9760 5057 9764
rect 5073 9820 5137 9824
rect 5073 9764 5077 9820
rect 5077 9764 5133 9820
rect 5133 9764 5137 9820
rect 5073 9760 5137 9764
rect 5153 9820 5217 9824
rect 5153 9764 5157 9820
rect 5157 9764 5213 9820
rect 5213 9764 5217 9820
rect 5153 9760 5217 9764
rect 5233 9820 5297 9824
rect 5233 9764 5237 9820
rect 5237 9764 5293 9820
rect 5293 9764 5297 9820
rect 5233 9760 5297 9764
rect 7247 9820 7311 9824
rect 7247 9764 7251 9820
rect 7251 9764 7307 9820
rect 7307 9764 7311 9820
rect 7247 9760 7311 9764
rect 7327 9820 7391 9824
rect 7327 9764 7331 9820
rect 7331 9764 7387 9820
rect 7387 9764 7391 9820
rect 7327 9760 7391 9764
rect 7407 9820 7471 9824
rect 7407 9764 7411 9820
rect 7411 9764 7467 9820
rect 7467 9764 7471 9820
rect 7407 9760 7471 9764
rect 7487 9820 7551 9824
rect 7487 9764 7491 9820
rect 7491 9764 7547 9820
rect 7547 9764 7551 9820
rect 7487 9760 7551 9764
rect 9501 9820 9565 9824
rect 9501 9764 9505 9820
rect 9505 9764 9561 9820
rect 9561 9764 9565 9820
rect 9501 9760 9565 9764
rect 9581 9820 9645 9824
rect 9581 9764 9585 9820
rect 9585 9764 9641 9820
rect 9641 9764 9645 9820
rect 9581 9760 9645 9764
rect 9661 9820 9725 9824
rect 9661 9764 9665 9820
rect 9665 9764 9721 9820
rect 9721 9764 9725 9820
rect 9661 9760 9725 9764
rect 9741 9820 9805 9824
rect 9741 9764 9745 9820
rect 9745 9764 9801 9820
rect 9801 9764 9805 9820
rect 9741 9760 9805 9764
rect 2079 9276 2143 9280
rect 2079 9220 2083 9276
rect 2083 9220 2139 9276
rect 2139 9220 2143 9276
rect 2079 9216 2143 9220
rect 2159 9276 2223 9280
rect 2159 9220 2163 9276
rect 2163 9220 2219 9276
rect 2219 9220 2223 9276
rect 2159 9216 2223 9220
rect 2239 9276 2303 9280
rect 2239 9220 2243 9276
rect 2243 9220 2299 9276
rect 2299 9220 2303 9276
rect 2239 9216 2303 9220
rect 2319 9276 2383 9280
rect 2319 9220 2323 9276
rect 2323 9220 2379 9276
rect 2379 9220 2383 9276
rect 2319 9216 2383 9220
rect 4333 9276 4397 9280
rect 4333 9220 4337 9276
rect 4337 9220 4393 9276
rect 4393 9220 4397 9276
rect 4333 9216 4397 9220
rect 4413 9276 4477 9280
rect 4413 9220 4417 9276
rect 4417 9220 4473 9276
rect 4473 9220 4477 9276
rect 4413 9216 4477 9220
rect 4493 9276 4557 9280
rect 4493 9220 4497 9276
rect 4497 9220 4553 9276
rect 4553 9220 4557 9276
rect 4493 9216 4557 9220
rect 4573 9276 4637 9280
rect 4573 9220 4577 9276
rect 4577 9220 4633 9276
rect 4633 9220 4637 9276
rect 4573 9216 4637 9220
rect 6587 9276 6651 9280
rect 6587 9220 6591 9276
rect 6591 9220 6647 9276
rect 6647 9220 6651 9276
rect 6587 9216 6651 9220
rect 6667 9276 6731 9280
rect 6667 9220 6671 9276
rect 6671 9220 6727 9276
rect 6727 9220 6731 9276
rect 6667 9216 6731 9220
rect 6747 9276 6811 9280
rect 6747 9220 6751 9276
rect 6751 9220 6807 9276
rect 6807 9220 6811 9276
rect 6747 9216 6811 9220
rect 6827 9276 6891 9280
rect 6827 9220 6831 9276
rect 6831 9220 6887 9276
rect 6887 9220 6891 9276
rect 6827 9216 6891 9220
rect 8841 9276 8905 9280
rect 8841 9220 8845 9276
rect 8845 9220 8901 9276
rect 8901 9220 8905 9276
rect 8841 9216 8905 9220
rect 8921 9276 8985 9280
rect 8921 9220 8925 9276
rect 8925 9220 8981 9276
rect 8981 9220 8985 9276
rect 8921 9216 8985 9220
rect 9001 9276 9065 9280
rect 9001 9220 9005 9276
rect 9005 9220 9061 9276
rect 9061 9220 9065 9276
rect 9001 9216 9065 9220
rect 9081 9276 9145 9280
rect 9081 9220 9085 9276
rect 9085 9220 9141 9276
rect 9141 9220 9145 9276
rect 9081 9216 9145 9220
rect 2739 8732 2803 8736
rect 2739 8676 2743 8732
rect 2743 8676 2799 8732
rect 2799 8676 2803 8732
rect 2739 8672 2803 8676
rect 2819 8732 2883 8736
rect 2819 8676 2823 8732
rect 2823 8676 2879 8732
rect 2879 8676 2883 8732
rect 2819 8672 2883 8676
rect 2899 8732 2963 8736
rect 2899 8676 2903 8732
rect 2903 8676 2959 8732
rect 2959 8676 2963 8732
rect 2899 8672 2963 8676
rect 2979 8732 3043 8736
rect 2979 8676 2983 8732
rect 2983 8676 3039 8732
rect 3039 8676 3043 8732
rect 2979 8672 3043 8676
rect 4993 8732 5057 8736
rect 4993 8676 4997 8732
rect 4997 8676 5053 8732
rect 5053 8676 5057 8732
rect 4993 8672 5057 8676
rect 5073 8732 5137 8736
rect 5073 8676 5077 8732
rect 5077 8676 5133 8732
rect 5133 8676 5137 8732
rect 5073 8672 5137 8676
rect 5153 8732 5217 8736
rect 5153 8676 5157 8732
rect 5157 8676 5213 8732
rect 5213 8676 5217 8732
rect 5153 8672 5217 8676
rect 5233 8732 5297 8736
rect 5233 8676 5237 8732
rect 5237 8676 5293 8732
rect 5293 8676 5297 8732
rect 5233 8672 5297 8676
rect 7247 8732 7311 8736
rect 7247 8676 7251 8732
rect 7251 8676 7307 8732
rect 7307 8676 7311 8732
rect 7247 8672 7311 8676
rect 7327 8732 7391 8736
rect 7327 8676 7331 8732
rect 7331 8676 7387 8732
rect 7387 8676 7391 8732
rect 7327 8672 7391 8676
rect 7407 8732 7471 8736
rect 7407 8676 7411 8732
rect 7411 8676 7467 8732
rect 7467 8676 7471 8732
rect 7407 8672 7471 8676
rect 7487 8732 7551 8736
rect 7487 8676 7491 8732
rect 7491 8676 7547 8732
rect 7547 8676 7551 8732
rect 7487 8672 7551 8676
rect 9501 8732 9565 8736
rect 9501 8676 9505 8732
rect 9505 8676 9561 8732
rect 9561 8676 9565 8732
rect 9501 8672 9565 8676
rect 9581 8732 9645 8736
rect 9581 8676 9585 8732
rect 9585 8676 9641 8732
rect 9641 8676 9645 8732
rect 9581 8672 9645 8676
rect 9661 8732 9725 8736
rect 9661 8676 9665 8732
rect 9665 8676 9721 8732
rect 9721 8676 9725 8732
rect 9661 8672 9725 8676
rect 9741 8732 9805 8736
rect 9741 8676 9745 8732
rect 9745 8676 9801 8732
rect 9801 8676 9805 8732
rect 9741 8672 9805 8676
rect 2079 8188 2143 8192
rect 2079 8132 2083 8188
rect 2083 8132 2139 8188
rect 2139 8132 2143 8188
rect 2079 8128 2143 8132
rect 2159 8188 2223 8192
rect 2159 8132 2163 8188
rect 2163 8132 2219 8188
rect 2219 8132 2223 8188
rect 2159 8128 2223 8132
rect 2239 8188 2303 8192
rect 2239 8132 2243 8188
rect 2243 8132 2299 8188
rect 2299 8132 2303 8188
rect 2239 8128 2303 8132
rect 2319 8188 2383 8192
rect 2319 8132 2323 8188
rect 2323 8132 2379 8188
rect 2379 8132 2383 8188
rect 2319 8128 2383 8132
rect 4333 8188 4397 8192
rect 4333 8132 4337 8188
rect 4337 8132 4393 8188
rect 4393 8132 4397 8188
rect 4333 8128 4397 8132
rect 4413 8188 4477 8192
rect 4413 8132 4417 8188
rect 4417 8132 4473 8188
rect 4473 8132 4477 8188
rect 4413 8128 4477 8132
rect 4493 8188 4557 8192
rect 4493 8132 4497 8188
rect 4497 8132 4553 8188
rect 4553 8132 4557 8188
rect 4493 8128 4557 8132
rect 4573 8188 4637 8192
rect 4573 8132 4577 8188
rect 4577 8132 4633 8188
rect 4633 8132 4637 8188
rect 4573 8128 4637 8132
rect 6587 8188 6651 8192
rect 6587 8132 6591 8188
rect 6591 8132 6647 8188
rect 6647 8132 6651 8188
rect 6587 8128 6651 8132
rect 6667 8188 6731 8192
rect 6667 8132 6671 8188
rect 6671 8132 6727 8188
rect 6727 8132 6731 8188
rect 6667 8128 6731 8132
rect 6747 8188 6811 8192
rect 6747 8132 6751 8188
rect 6751 8132 6807 8188
rect 6807 8132 6811 8188
rect 6747 8128 6811 8132
rect 6827 8188 6891 8192
rect 6827 8132 6831 8188
rect 6831 8132 6887 8188
rect 6887 8132 6891 8188
rect 6827 8128 6891 8132
rect 8841 8188 8905 8192
rect 8841 8132 8845 8188
rect 8845 8132 8901 8188
rect 8901 8132 8905 8188
rect 8841 8128 8905 8132
rect 8921 8188 8985 8192
rect 8921 8132 8925 8188
rect 8925 8132 8981 8188
rect 8981 8132 8985 8188
rect 8921 8128 8985 8132
rect 9001 8188 9065 8192
rect 9001 8132 9005 8188
rect 9005 8132 9061 8188
rect 9061 8132 9065 8188
rect 9001 8128 9065 8132
rect 9081 8188 9145 8192
rect 9081 8132 9085 8188
rect 9085 8132 9141 8188
rect 9141 8132 9145 8188
rect 9081 8128 9145 8132
rect 2739 7644 2803 7648
rect 2739 7588 2743 7644
rect 2743 7588 2799 7644
rect 2799 7588 2803 7644
rect 2739 7584 2803 7588
rect 2819 7644 2883 7648
rect 2819 7588 2823 7644
rect 2823 7588 2879 7644
rect 2879 7588 2883 7644
rect 2819 7584 2883 7588
rect 2899 7644 2963 7648
rect 2899 7588 2903 7644
rect 2903 7588 2959 7644
rect 2959 7588 2963 7644
rect 2899 7584 2963 7588
rect 2979 7644 3043 7648
rect 2979 7588 2983 7644
rect 2983 7588 3039 7644
rect 3039 7588 3043 7644
rect 2979 7584 3043 7588
rect 4993 7644 5057 7648
rect 4993 7588 4997 7644
rect 4997 7588 5053 7644
rect 5053 7588 5057 7644
rect 4993 7584 5057 7588
rect 5073 7644 5137 7648
rect 5073 7588 5077 7644
rect 5077 7588 5133 7644
rect 5133 7588 5137 7644
rect 5073 7584 5137 7588
rect 5153 7644 5217 7648
rect 5153 7588 5157 7644
rect 5157 7588 5213 7644
rect 5213 7588 5217 7644
rect 5153 7584 5217 7588
rect 5233 7644 5297 7648
rect 5233 7588 5237 7644
rect 5237 7588 5293 7644
rect 5293 7588 5297 7644
rect 5233 7584 5297 7588
rect 7247 7644 7311 7648
rect 7247 7588 7251 7644
rect 7251 7588 7307 7644
rect 7307 7588 7311 7644
rect 7247 7584 7311 7588
rect 7327 7644 7391 7648
rect 7327 7588 7331 7644
rect 7331 7588 7387 7644
rect 7387 7588 7391 7644
rect 7327 7584 7391 7588
rect 7407 7644 7471 7648
rect 7407 7588 7411 7644
rect 7411 7588 7467 7644
rect 7467 7588 7471 7644
rect 7407 7584 7471 7588
rect 7487 7644 7551 7648
rect 7487 7588 7491 7644
rect 7491 7588 7547 7644
rect 7547 7588 7551 7644
rect 7487 7584 7551 7588
rect 9501 7644 9565 7648
rect 9501 7588 9505 7644
rect 9505 7588 9561 7644
rect 9561 7588 9565 7644
rect 9501 7584 9565 7588
rect 9581 7644 9645 7648
rect 9581 7588 9585 7644
rect 9585 7588 9641 7644
rect 9641 7588 9645 7644
rect 9581 7584 9645 7588
rect 9661 7644 9725 7648
rect 9661 7588 9665 7644
rect 9665 7588 9721 7644
rect 9721 7588 9725 7644
rect 9661 7584 9725 7588
rect 9741 7644 9805 7648
rect 9741 7588 9745 7644
rect 9745 7588 9801 7644
rect 9801 7588 9805 7644
rect 9741 7584 9805 7588
rect 2079 7100 2143 7104
rect 2079 7044 2083 7100
rect 2083 7044 2139 7100
rect 2139 7044 2143 7100
rect 2079 7040 2143 7044
rect 2159 7100 2223 7104
rect 2159 7044 2163 7100
rect 2163 7044 2219 7100
rect 2219 7044 2223 7100
rect 2159 7040 2223 7044
rect 2239 7100 2303 7104
rect 2239 7044 2243 7100
rect 2243 7044 2299 7100
rect 2299 7044 2303 7100
rect 2239 7040 2303 7044
rect 2319 7100 2383 7104
rect 2319 7044 2323 7100
rect 2323 7044 2379 7100
rect 2379 7044 2383 7100
rect 2319 7040 2383 7044
rect 4333 7100 4397 7104
rect 4333 7044 4337 7100
rect 4337 7044 4393 7100
rect 4393 7044 4397 7100
rect 4333 7040 4397 7044
rect 4413 7100 4477 7104
rect 4413 7044 4417 7100
rect 4417 7044 4473 7100
rect 4473 7044 4477 7100
rect 4413 7040 4477 7044
rect 4493 7100 4557 7104
rect 4493 7044 4497 7100
rect 4497 7044 4553 7100
rect 4553 7044 4557 7100
rect 4493 7040 4557 7044
rect 4573 7100 4637 7104
rect 4573 7044 4577 7100
rect 4577 7044 4633 7100
rect 4633 7044 4637 7100
rect 4573 7040 4637 7044
rect 6587 7100 6651 7104
rect 6587 7044 6591 7100
rect 6591 7044 6647 7100
rect 6647 7044 6651 7100
rect 6587 7040 6651 7044
rect 6667 7100 6731 7104
rect 6667 7044 6671 7100
rect 6671 7044 6727 7100
rect 6727 7044 6731 7100
rect 6667 7040 6731 7044
rect 6747 7100 6811 7104
rect 6747 7044 6751 7100
rect 6751 7044 6807 7100
rect 6807 7044 6811 7100
rect 6747 7040 6811 7044
rect 6827 7100 6891 7104
rect 6827 7044 6831 7100
rect 6831 7044 6887 7100
rect 6887 7044 6891 7100
rect 6827 7040 6891 7044
rect 8841 7100 8905 7104
rect 8841 7044 8845 7100
rect 8845 7044 8901 7100
rect 8901 7044 8905 7100
rect 8841 7040 8905 7044
rect 8921 7100 8985 7104
rect 8921 7044 8925 7100
rect 8925 7044 8981 7100
rect 8981 7044 8985 7100
rect 8921 7040 8985 7044
rect 9001 7100 9065 7104
rect 9001 7044 9005 7100
rect 9005 7044 9061 7100
rect 9061 7044 9065 7100
rect 9001 7040 9065 7044
rect 9081 7100 9145 7104
rect 9081 7044 9085 7100
rect 9085 7044 9141 7100
rect 9141 7044 9145 7100
rect 9081 7040 9145 7044
rect 4108 7032 4172 7036
rect 4108 6976 4158 7032
rect 4158 6976 4172 7032
rect 4108 6972 4172 6976
rect 2739 6556 2803 6560
rect 2739 6500 2743 6556
rect 2743 6500 2799 6556
rect 2799 6500 2803 6556
rect 2739 6496 2803 6500
rect 2819 6556 2883 6560
rect 2819 6500 2823 6556
rect 2823 6500 2879 6556
rect 2879 6500 2883 6556
rect 2819 6496 2883 6500
rect 2899 6556 2963 6560
rect 2899 6500 2903 6556
rect 2903 6500 2959 6556
rect 2959 6500 2963 6556
rect 2899 6496 2963 6500
rect 2979 6556 3043 6560
rect 2979 6500 2983 6556
rect 2983 6500 3039 6556
rect 3039 6500 3043 6556
rect 2979 6496 3043 6500
rect 4993 6556 5057 6560
rect 4993 6500 4997 6556
rect 4997 6500 5053 6556
rect 5053 6500 5057 6556
rect 4993 6496 5057 6500
rect 5073 6556 5137 6560
rect 5073 6500 5077 6556
rect 5077 6500 5133 6556
rect 5133 6500 5137 6556
rect 5073 6496 5137 6500
rect 5153 6556 5217 6560
rect 5153 6500 5157 6556
rect 5157 6500 5213 6556
rect 5213 6500 5217 6556
rect 5153 6496 5217 6500
rect 5233 6556 5297 6560
rect 5233 6500 5237 6556
rect 5237 6500 5293 6556
rect 5293 6500 5297 6556
rect 5233 6496 5297 6500
rect 7247 6556 7311 6560
rect 7247 6500 7251 6556
rect 7251 6500 7307 6556
rect 7307 6500 7311 6556
rect 7247 6496 7311 6500
rect 7327 6556 7391 6560
rect 7327 6500 7331 6556
rect 7331 6500 7387 6556
rect 7387 6500 7391 6556
rect 7327 6496 7391 6500
rect 7407 6556 7471 6560
rect 7407 6500 7411 6556
rect 7411 6500 7467 6556
rect 7467 6500 7471 6556
rect 7407 6496 7471 6500
rect 7487 6556 7551 6560
rect 7487 6500 7491 6556
rect 7491 6500 7547 6556
rect 7547 6500 7551 6556
rect 7487 6496 7551 6500
rect 9501 6556 9565 6560
rect 9501 6500 9505 6556
rect 9505 6500 9561 6556
rect 9561 6500 9565 6556
rect 9501 6496 9565 6500
rect 9581 6556 9645 6560
rect 9581 6500 9585 6556
rect 9585 6500 9641 6556
rect 9641 6500 9645 6556
rect 9581 6496 9645 6500
rect 9661 6556 9725 6560
rect 9661 6500 9665 6556
rect 9665 6500 9721 6556
rect 9721 6500 9725 6556
rect 9661 6496 9725 6500
rect 9741 6556 9805 6560
rect 9741 6500 9745 6556
rect 9745 6500 9801 6556
rect 9801 6500 9805 6556
rect 9741 6496 9805 6500
rect 2079 6012 2143 6016
rect 2079 5956 2083 6012
rect 2083 5956 2139 6012
rect 2139 5956 2143 6012
rect 2079 5952 2143 5956
rect 2159 6012 2223 6016
rect 2159 5956 2163 6012
rect 2163 5956 2219 6012
rect 2219 5956 2223 6012
rect 2159 5952 2223 5956
rect 2239 6012 2303 6016
rect 2239 5956 2243 6012
rect 2243 5956 2299 6012
rect 2299 5956 2303 6012
rect 2239 5952 2303 5956
rect 2319 6012 2383 6016
rect 2319 5956 2323 6012
rect 2323 5956 2379 6012
rect 2379 5956 2383 6012
rect 2319 5952 2383 5956
rect 4333 6012 4397 6016
rect 4333 5956 4337 6012
rect 4337 5956 4393 6012
rect 4393 5956 4397 6012
rect 4333 5952 4397 5956
rect 4413 6012 4477 6016
rect 4413 5956 4417 6012
rect 4417 5956 4473 6012
rect 4473 5956 4477 6012
rect 4413 5952 4477 5956
rect 4493 6012 4557 6016
rect 4493 5956 4497 6012
rect 4497 5956 4553 6012
rect 4553 5956 4557 6012
rect 4493 5952 4557 5956
rect 4573 6012 4637 6016
rect 4573 5956 4577 6012
rect 4577 5956 4633 6012
rect 4633 5956 4637 6012
rect 4573 5952 4637 5956
rect 6587 6012 6651 6016
rect 6587 5956 6591 6012
rect 6591 5956 6647 6012
rect 6647 5956 6651 6012
rect 6587 5952 6651 5956
rect 6667 6012 6731 6016
rect 6667 5956 6671 6012
rect 6671 5956 6727 6012
rect 6727 5956 6731 6012
rect 6667 5952 6731 5956
rect 6747 6012 6811 6016
rect 6747 5956 6751 6012
rect 6751 5956 6807 6012
rect 6807 5956 6811 6012
rect 6747 5952 6811 5956
rect 6827 6012 6891 6016
rect 6827 5956 6831 6012
rect 6831 5956 6887 6012
rect 6887 5956 6891 6012
rect 6827 5952 6891 5956
rect 8841 6012 8905 6016
rect 8841 5956 8845 6012
rect 8845 5956 8901 6012
rect 8901 5956 8905 6012
rect 8841 5952 8905 5956
rect 8921 6012 8985 6016
rect 8921 5956 8925 6012
rect 8925 5956 8981 6012
rect 8981 5956 8985 6012
rect 8921 5952 8985 5956
rect 9001 6012 9065 6016
rect 9001 5956 9005 6012
rect 9005 5956 9061 6012
rect 9061 5956 9065 6012
rect 9001 5952 9065 5956
rect 9081 6012 9145 6016
rect 9081 5956 9085 6012
rect 9085 5956 9141 6012
rect 9141 5956 9145 6012
rect 9081 5952 9145 5956
rect 2739 5468 2803 5472
rect 2739 5412 2743 5468
rect 2743 5412 2799 5468
rect 2799 5412 2803 5468
rect 2739 5408 2803 5412
rect 2819 5468 2883 5472
rect 2819 5412 2823 5468
rect 2823 5412 2879 5468
rect 2879 5412 2883 5468
rect 2819 5408 2883 5412
rect 2899 5468 2963 5472
rect 2899 5412 2903 5468
rect 2903 5412 2959 5468
rect 2959 5412 2963 5468
rect 2899 5408 2963 5412
rect 2979 5468 3043 5472
rect 2979 5412 2983 5468
rect 2983 5412 3039 5468
rect 3039 5412 3043 5468
rect 2979 5408 3043 5412
rect 4993 5468 5057 5472
rect 4993 5412 4997 5468
rect 4997 5412 5053 5468
rect 5053 5412 5057 5468
rect 4993 5408 5057 5412
rect 5073 5468 5137 5472
rect 5073 5412 5077 5468
rect 5077 5412 5133 5468
rect 5133 5412 5137 5468
rect 5073 5408 5137 5412
rect 5153 5468 5217 5472
rect 5153 5412 5157 5468
rect 5157 5412 5213 5468
rect 5213 5412 5217 5468
rect 5153 5408 5217 5412
rect 5233 5468 5297 5472
rect 5233 5412 5237 5468
rect 5237 5412 5293 5468
rect 5293 5412 5297 5468
rect 5233 5408 5297 5412
rect 7247 5468 7311 5472
rect 7247 5412 7251 5468
rect 7251 5412 7307 5468
rect 7307 5412 7311 5468
rect 7247 5408 7311 5412
rect 7327 5468 7391 5472
rect 7327 5412 7331 5468
rect 7331 5412 7387 5468
rect 7387 5412 7391 5468
rect 7327 5408 7391 5412
rect 7407 5468 7471 5472
rect 7407 5412 7411 5468
rect 7411 5412 7467 5468
rect 7467 5412 7471 5468
rect 7407 5408 7471 5412
rect 7487 5468 7551 5472
rect 7487 5412 7491 5468
rect 7491 5412 7547 5468
rect 7547 5412 7551 5468
rect 7487 5408 7551 5412
rect 9501 5468 9565 5472
rect 9501 5412 9505 5468
rect 9505 5412 9561 5468
rect 9561 5412 9565 5468
rect 9501 5408 9565 5412
rect 9581 5468 9645 5472
rect 9581 5412 9585 5468
rect 9585 5412 9641 5468
rect 9641 5412 9645 5468
rect 9581 5408 9645 5412
rect 9661 5468 9725 5472
rect 9661 5412 9665 5468
rect 9665 5412 9721 5468
rect 9721 5412 9725 5468
rect 9661 5408 9725 5412
rect 9741 5468 9805 5472
rect 9741 5412 9745 5468
rect 9745 5412 9801 5468
rect 9801 5412 9805 5468
rect 9741 5408 9805 5412
rect 2079 4924 2143 4928
rect 2079 4868 2083 4924
rect 2083 4868 2139 4924
rect 2139 4868 2143 4924
rect 2079 4864 2143 4868
rect 2159 4924 2223 4928
rect 2159 4868 2163 4924
rect 2163 4868 2219 4924
rect 2219 4868 2223 4924
rect 2159 4864 2223 4868
rect 2239 4924 2303 4928
rect 2239 4868 2243 4924
rect 2243 4868 2299 4924
rect 2299 4868 2303 4924
rect 2239 4864 2303 4868
rect 2319 4924 2383 4928
rect 2319 4868 2323 4924
rect 2323 4868 2379 4924
rect 2379 4868 2383 4924
rect 2319 4864 2383 4868
rect 4333 4924 4397 4928
rect 4333 4868 4337 4924
rect 4337 4868 4393 4924
rect 4393 4868 4397 4924
rect 4333 4864 4397 4868
rect 4413 4924 4477 4928
rect 4413 4868 4417 4924
rect 4417 4868 4473 4924
rect 4473 4868 4477 4924
rect 4413 4864 4477 4868
rect 4493 4924 4557 4928
rect 4493 4868 4497 4924
rect 4497 4868 4553 4924
rect 4553 4868 4557 4924
rect 4493 4864 4557 4868
rect 4573 4924 4637 4928
rect 4573 4868 4577 4924
rect 4577 4868 4633 4924
rect 4633 4868 4637 4924
rect 4573 4864 4637 4868
rect 6587 4924 6651 4928
rect 6587 4868 6591 4924
rect 6591 4868 6647 4924
rect 6647 4868 6651 4924
rect 6587 4864 6651 4868
rect 6667 4924 6731 4928
rect 6667 4868 6671 4924
rect 6671 4868 6727 4924
rect 6727 4868 6731 4924
rect 6667 4864 6731 4868
rect 6747 4924 6811 4928
rect 6747 4868 6751 4924
rect 6751 4868 6807 4924
rect 6807 4868 6811 4924
rect 6747 4864 6811 4868
rect 6827 4924 6891 4928
rect 6827 4868 6831 4924
rect 6831 4868 6887 4924
rect 6887 4868 6891 4924
rect 6827 4864 6891 4868
rect 8841 4924 8905 4928
rect 8841 4868 8845 4924
rect 8845 4868 8901 4924
rect 8901 4868 8905 4924
rect 8841 4864 8905 4868
rect 8921 4924 8985 4928
rect 8921 4868 8925 4924
rect 8925 4868 8981 4924
rect 8981 4868 8985 4924
rect 8921 4864 8985 4868
rect 9001 4924 9065 4928
rect 9001 4868 9005 4924
rect 9005 4868 9061 4924
rect 9061 4868 9065 4924
rect 9001 4864 9065 4868
rect 9081 4924 9145 4928
rect 9081 4868 9085 4924
rect 9085 4868 9141 4924
rect 9141 4868 9145 4924
rect 9081 4864 9145 4868
rect 2739 4380 2803 4384
rect 2739 4324 2743 4380
rect 2743 4324 2799 4380
rect 2799 4324 2803 4380
rect 2739 4320 2803 4324
rect 2819 4380 2883 4384
rect 2819 4324 2823 4380
rect 2823 4324 2879 4380
rect 2879 4324 2883 4380
rect 2819 4320 2883 4324
rect 2899 4380 2963 4384
rect 2899 4324 2903 4380
rect 2903 4324 2959 4380
rect 2959 4324 2963 4380
rect 2899 4320 2963 4324
rect 2979 4380 3043 4384
rect 2979 4324 2983 4380
rect 2983 4324 3039 4380
rect 3039 4324 3043 4380
rect 2979 4320 3043 4324
rect 4993 4380 5057 4384
rect 4993 4324 4997 4380
rect 4997 4324 5053 4380
rect 5053 4324 5057 4380
rect 4993 4320 5057 4324
rect 5073 4380 5137 4384
rect 5073 4324 5077 4380
rect 5077 4324 5133 4380
rect 5133 4324 5137 4380
rect 5073 4320 5137 4324
rect 5153 4380 5217 4384
rect 5153 4324 5157 4380
rect 5157 4324 5213 4380
rect 5213 4324 5217 4380
rect 5153 4320 5217 4324
rect 5233 4380 5297 4384
rect 5233 4324 5237 4380
rect 5237 4324 5293 4380
rect 5293 4324 5297 4380
rect 5233 4320 5297 4324
rect 7247 4380 7311 4384
rect 7247 4324 7251 4380
rect 7251 4324 7307 4380
rect 7307 4324 7311 4380
rect 7247 4320 7311 4324
rect 7327 4380 7391 4384
rect 7327 4324 7331 4380
rect 7331 4324 7387 4380
rect 7387 4324 7391 4380
rect 7327 4320 7391 4324
rect 7407 4380 7471 4384
rect 7407 4324 7411 4380
rect 7411 4324 7467 4380
rect 7467 4324 7471 4380
rect 7407 4320 7471 4324
rect 7487 4380 7551 4384
rect 7487 4324 7491 4380
rect 7491 4324 7547 4380
rect 7547 4324 7551 4380
rect 7487 4320 7551 4324
rect 9501 4380 9565 4384
rect 9501 4324 9505 4380
rect 9505 4324 9561 4380
rect 9561 4324 9565 4380
rect 9501 4320 9565 4324
rect 9581 4380 9645 4384
rect 9581 4324 9585 4380
rect 9585 4324 9641 4380
rect 9641 4324 9645 4380
rect 9581 4320 9645 4324
rect 9661 4380 9725 4384
rect 9661 4324 9665 4380
rect 9665 4324 9721 4380
rect 9721 4324 9725 4380
rect 9661 4320 9725 4324
rect 9741 4380 9805 4384
rect 9741 4324 9745 4380
rect 9745 4324 9801 4380
rect 9801 4324 9805 4380
rect 9741 4320 9805 4324
rect 4108 3980 4172 4044
rect 2079 3836 2143 3840
rect 2079 3780 2083 3836
rect 2083 3780 2139 3836
rect 2139 3780 2143 3836
rect 2079 3776 2143 3780
rect 2159 3836 2223 3840
rect 2159 3780 2163 3836
rect 2163 3780 2219 3836
rect 2219 3780 2223 3836
rect 2159 3776 2223 3780
rect 2239 3836 2303 3840
rect 2239 3780 2243 3836
rect 2243 3780 2299 3836
rect 2299 3780 2303 3836
rect 2239 3776 2303 3780
rect 2319 3836 2383 3840
rect 2319 3780 2323 3836
rect 2323 3780 2379 3836
rect 2379 3780 2383 3836
rect 2319 3776 2383 3780
rect 4333 3836 4397 3840
rect 4333 3780 4337 3836
rect 4337 3780 4393 3836
rect 4393 3780 4397 3836
rect 4333 3776 4397 3780
rect 4413 3836 4477 3840
rect 4413 3780 4417 3836
rect 4417 3780 4473 3836
rect 4473 3780 4477 3836
rect 4413 3776 4477 3780
rect 4493 3836 4557 3840
rect 4493 3780 4497 3836
rect 4497 3780 4553 3836
rect 4553 3780 4557 3836
rect 4493 3776 4557 3780
rect 4573 3836 4637 3840
rect 4573 3780 4577 3836
rect 4577 3780 4633 3836
rect 4633 3780 4637 3836
rect 4573 3776 4637 3780
rect 6587 3836 6651 3840
rect 6587 3780 6591 3836
rect 6591 3780 6647 3836
rect 6647 3780 6651 3836
rect 6587 3776 6651 3780
rect 6667 3836 6731 3840
rect 6667 3780 6671 3836
rect 6671 3780 6727 3836
rect 6727 3780 6731 3836
rect 6667 3776 6731 3780
rect 6747 3836 6811 3840
rect 6747 3780 6751 3836
rect 6751 3780 6807 3836
rect 6807 3780 6811 3836
rect 6747 3776 6811 3780
rect 6827 3836 6891 3840
rect 6827 3780 6831 3836
rect 6831 3780 6887 3836
rect 6887 3780 6891 3836
rect 6827 3776 6891 3780
rect 8841 3836 8905 3840
rect 8841 3780 8845 3836
rect 8845 3780 8901 3836
rect 8901 3780 8905 3836
rect 8841 3776 8905 3780
rect 8921 3836 8985 3840
rect 8921 3780 8925 3836
rect 8925 3780 8981 3836
rect 8981 3780 8985 3836
rect 8921 3776 8985 3780
rect 9001 3836 9065 3840
rect 9001 3780 9005 3836
rect 9005 3780 9061 3836
rect 9061 3780 9065 3836
rect 9001 3776 9065 3780
rect 9081 3836 9145 3840
rect 9081 3780 9085 3836
rect 9085 3780 9141 3836
rect 9141 3780 9145 3836
rect 9081 3776 9145 3780
rect 2739 3292 2803 3296
rect 2739 3236 2743 3292
rect 2743 3236 2799 3292
rect 2799 3236 2803 3292
rect 2739 3232 2803 3236
rect 2819 3292 2883 3296
rect 2819 3236 2823 3292
rect 2823 3236 2879 3292
rect 2879 3236 2883 3292
rect 2819 3232 2883 3236
rect 2899 3292 2963 3296
rect 2899 3236 2903 3292
rect 2903 3236 2959 3292
rect 2959 3236 2963 3292
rect 2899 3232 2963 3236
rect 2979 3292 3043 3296
rect 2979 3236 2983 3292
rect 2983 3236 3039 3292
rect 3039 3236 3043 3292
rect 2979 3232 3043 3236
rect 4993 3292 5057 3296
rect 4993 3236 4997 3292
rect 4997 3236 5053 3292
rect 5053 3236 5057 3292
rect 4993 3232 5057 3236
rect 5073 3292 5137 3296
rect 5073 3236 5077 3292
rect 5077 3236 5133 3292
rect 5133 3236 5137 3292
rect 5073 3232 5137 3236
rect 5153 3292 5217 3296
rect 5153 3236 5157 3292
rect 5157 3236 5213 3292
rect 5213 3236 5217 3292
rect 5153 3232 5217 3236
rect 5233 3292 5297 3296
rect 5233 3236 5237 3292
rect 5237 3236 5293 3292
rect 5293 3236 5297 3292
rect 5233 3232 5297 3236
rect 7247 3292 7311 3296
rect 7247 3236 7251 3292
rect 7251 3236 7307 3292
rect 7307 3236 7311 3292
rect 7247 3232 7311 3236
rect 7327 3292 7391 3296
rect 7327 3236 7331 3292
rect 7331 3236 7387 3292
rect 7387 3236 7391 3292
rect 7327 3232 7391 3236
rect 7407 3292 7471 3296
rect 7407 3236 7411 3292
rect 7411 3236 7467 3292
rect 7467 3236 7471 3292
rect 7407 3232 7471 3236
rect 7487 3292 7551 3296
rect 7487 3236 7491 3292
rect 7491 3236 7547 3292
rect 7547 3236 7551 3292
rect 7487 3232 7551 3236
rect 9501 3292 9565 3296
rect 9501 3236 9505 3292
rect 9505 3236 9561 3292
rect 9561 3236 9565 3292
rect 9501 3232 9565 3236
rect 9581 3292 9645 3296
rect 9581 3236 9585 3292
rect 9585 3236 9641 3292
rect 9641 3236 9645 3292
rect 9581 3232 9645 3236
rect 9661 3292 9725 3296
rect 9661 3236 9665 3292
rect 9665 3236 9721 3292
rect 9721 3236 9725 3292
rect 9661 3232 9725 3236
rect 9741 3292 9805 3296
rect 9741 3236 9745 3292
rect 9745 3236 9801 3292
rect 9801 3236 9805 3292
rect 9741 3232 9805 3236
rect 2079 2748 2143 2752
rect 2079 2692 2083 2748
rect 2083 2692 2139 2748
rect 2139 2692 2143 2748
rect 2079 2688 2143 2692
rect 2159 2748 2223 2752
rect 2159 2692 2163 2748
rect 2163 2692 2219 2748
rect 2219 2692 2223 2748
rect 2159 2688 2223 2692
rect 2239 2748 2303 2752
rect 2239 2692 2243 2748
rect 2243 2692 2299 2748
rect 2299 2692 2303 2748
rect 2239 2688 2303 2692
rect 2319 2748 2383 2752
rect 2319 2692 2323 2748
rect 2323 2692 2379 2748
rect 2379 2692 2383 2748
rect 2319 2688 2383 2692
rect 4333 2748 4397 2752
rect 4333 2692 4337 2748
rect 4337 2692 4393 2748
rect 4393 2692 4397 2748
rect 4333 2688 4397 2692
rect 4413 2748 4477 2752
rect 4413 2692 4417 2748
rect 4417 2692 4473 2748
rect 4473 2692 4477 2748
rect 4413 2688 4477 2692
rect 4493 2748 4557 2752
rect 4493 2692 4497 2748
rect 4497 2692 4553 2748
rect 4553 2692 4557 2748
rect 4493 2688 4557 2692
rect 4573 2748 4637 2752
rect 4573 2692 4577 2748
rect 4577 2692 4633 2748
rect 4633 2692 4637 2748
rect 4573 2688 4637 2692
rect 6587 2748 6651 2752
rect 6587 2692 6591 2748
rect 6591 2692 6647 2748
rect 6647 2692 6651 2748
rect 6587 2688 6651 2692
rect 6667 2748 6731 2752
rect 6667 2692 6671 2748
rect 6671 2692 6727 2748
rect 6727 2692 6731 2748
rect 6667 2688 6731 2692
rect 6747 2748 6811 2752
rect 6747 2692 6751 2748
rect 6751 2692 6807 2748
rect 6807 2692 6811 2748
rect 6747 2688 6811 2692
rect 6827 2748 6891 2752
rect 6827 2692 6831 2748
rect 6831 2692 6887 2748
rect 6887 2692 6891 2748
rect 6827 2688 6891 2692
rect 8841 2748 8905 2752
rect 8841 2692 8845 2748
rect 8845 2692 8901 2748
rect 8901 2692 8905 2748
rect 8841 2688 8905 2692
rect 8921 2748 8985 2752
rect 8921 2692 8925 2748
rect 8925 2692 8981 2748
rect 8981 2692 8985 2748
rect 8921 2688 8985 2692
rect 9001 2748 9065 2752
rect 9001 2692 9005 2748
rect 9005 2692 9061 2748
rect 9061 2692 9065 2748
rect 9001 2688 9065 2692
rect 9081 2748 9145 2752
rect 9081 2692 9085 2748
rect 9085 2692 9141 2748
rect 9141 2692 9145 2748
rect 9081 2688 9145 2692
rect 2739 2204 2803 2208
rect 2739 2148 2743 2204
rect 2743 2148 2799 2204
rect 2799 2148 2803 2204
rect 2739 2144 2803 2148
rect 2819 2204 2883 2208
rect 2819 2148 2823 2204
rect 2823 2148 2879 2204
rect 2879 2148 2883 2204
rect 2819 2144 2883 2148
rect 2899 2204 2963 2208
rect 2899 2148 2903 2204
rect 2903 2148 2959 2204
rect 2959 2148 2963 2204
rect 2899 2144 2963 2148
rect 2979 2204 3043 2208
rect 2979 2148 2983 2204
rect 2983 2148 3039 2204
rect 3039 2148 3043 2204
rect 2979 2144 3043 2148
rect 4993 2204 5057 2208
rect 4993 2148 4997 2204
rect 4997 2148 5053 2204
rect 5053 2148 5057 2204
rect 4993 2144 5057 2148
rect 5073 2204 5137 2208
rect 5073 2148 5077 2204
rect 5077 2148 5133 2204
rect 5133 2148 5137 2204
rect 5073 2144 5137 2148
rect 5153 2204 5217 2208
rect 5153 2148 5157 2204
rect 5157 2148 5213 2204
rect 5213 2148 5217 2204
rect 5153 2144 5217 2148
rect 5233 2204 5297 2208
rect 5233 2148 5237 2204
rect 5237 2148 5293 2204
rect 5293 2148 5297 2204
rect 5233 2144 5297 2148
rect 7247 2204 7311 2208
rect 7247 2148 7251 2204
rect 7251 2148 7307 2204
rect 7307 2148 7311 2204
rect 7247 2144 7311 2148
rect 7327 2204 7391 2208
rect 7327 2148 7331 2204
rect 7331 2148 7387 2204
rect 7387 2148 7391 2204
rect 7327 2144 7391 2148
rect 7407 2204 7471 2208
rect 7407 2148 7411 2204
rect 7411 2148 7467 2204
rect 7467 2148 7471 2204
rect 7407 2144 7471 2148
rect 7487 2204 7551 2208
rect 7487 2148 7491 2204
rect 7491 2148 7547 2204
rect 7547 2148 7551 2204
rect 7487 2144 7551 2148
rect 9501 2204 9565 2208
rect 9501 2148 9505 2204
rect 9505 2148 9561 2204
rect 9561 2148 9565 2204
rect 9501 2144 9565 2148
rect 9581 2204 9645 2208
rect 9581 2148 9585 2204
rect 9585 2148 9641 2204
rect 9641 2148 9645 2204
rect 9581 2144 9645 2148
rect 9661 2204 9725 2208
rect 9661 2148 9665 2204
rect 9665 2148 9721 2204
rect 9721 2148 9725 2204
rect 9661 2144 9725 2148
rect 9741 2204 9805 2208
rect 9741 2148 9745 2204
rect 9745 2148 9801 2204
rect 9801 2148 9805 2204
rect 9741 2144 9805 2148
<< metal4 >>
rect 2071 10368 2391 10928
rect 2071 10304 2079 10368
rect 2143 10304 2159 10368
rect 2223 10304 2239 10368
rect 2303 10304 2319 10368
rect 2383 10304 2391 10368
rect 2071 9906 2391 10304
rect 2071 9670 2113 9906
rect 2349 9670 2391 9906
rect 2071 9280 2391 9670
rect 2071 9216 2079 9280
rect 2143 9216 2159 9280
rect 2223 9216 2239 9280
rect 2303 9216 2319 9280
rect 2383 9216 2391 9280
rect 2071 8192 2391 9216
rect 2071 8128 2079 8192
rect 2143 8128 2159 8192
rect 2223 8128 2239 8192
rect 2303 8128 2319 8192
rect 2383 8128 2391 8192
rect 2071 7731 2391 8128
rect 2071 7495 2113 7731
rect 2349 7495 2391 7731
rect 2071 7104 2391 7495
rect 2071 7040 2079 7104
rect 2143 7040 2159 7104
rect 2223 7040 2239 7104
rect 2303 7040 2319 7104
rect 2383 7040 2391 7104
rect 2071 6016 2391 7040
rect 2071 5952 2079 6016
rect 2143 5952 2159 6016
rect 2223 5952 2239 6016
rect 2303 5952 2319 6016
rect 2383 5952 2391 6016
rect 2071 5556 2391 5952
rect 2071 5320 2113 5556
rect 2349 5320 2391 5556
rect 2071 4928 2391 5320
rect 2071 4864 2079 4928
rect 2143 4864 2159 4928
rect 2223 4864 2239 4928
rect 2303 4864 2319 4928
rect 2383 4864 2391 4928
rect 2071 3840 2391 4864
rect 2071 3776 2079 3840
rect 2143 3776 2159 3840
rect 2223 3776 2239 3840
rect 2303 3776 2319 3840
rect 2383 3776 2391 3840
rect 2071 3381 2391 3776
rect 2071 3145 2113 3381
rect 2349 3145 2391 3381
rect 2071 2752 2391 3145
rect 2071 2688 2079 2752
rect 2143 2688 2159 2752
rect 2223 2688 2239 2752
rect 2303 2688 2319 2752
rect 2383 2688 2391 2752
rect 2071 2128 2391 2688
rect 2731 10912 3051 10928
rect 2731 10848 2739 10912
rect 2803 10848 2819 10912
rect 2883 10848 2899 10912
rect 2963 10848 2979 10912
rect 3043 10848 3051 10912
rect 2731 10566 3051 10848
rect 2731 10330 2773 10566
rect 3009 10330 3051 10566
rect 2731 9824 3051 10330
rect 2731 9760 2739 9824
rect 2803 9760 2819 9824
rect 2883 9760 2899 9824
rect 2963 9760 2979 9824
rect 3043 9760 3051 9824
rect 2731 8736 3051 9760
rect 2731 8672 2739 8736
rect 2803 8672 2819 8736
rect 2883 8672 2899 8736
rect 2963 8672 2979 8736
rect 3043 8672 3051 8736
rect 2731 8391 3051 8672
rect 2731 8155 2773 8391
rect 3009 8155 3051 8391
rect 2731 7648 3051 8155
rect 2731 7584 2739 7648
rect 2803 7584 2819 7648
rect 2883 7584 2899 7648
rect 2963 7584 2979 7648
rect 3043 7584 3051 7648
rect 2731 6560 3051 7584
rect 4325 10368 4645 10928
rect 4325 10304 4333 10368
rect 4397 10304 4413 10368
rect 4477 10304 4493 10368
rect 4557 10304 4573 10368
rect 4637 10304 4645 10368
rect 4325 9906 4645 10304
rect 4325 9670 4367 9906
rect 4603 9670 4645 9906
rect 4325 9280 4645 9670
rect 4325 9216 4333 9280
rect 4397 9216 4413 9280
rect 4477 9216 4493 9280
rect 4557 9216 4573 9280
rect 4637 9216 4645 9280
rect 4325 8192 4645 9216
rect 4325 8128 4333 8192
rect 4397 8128 4413 8192
rect 4477 8128 4493 8192
rect 4557 8128 4573 8192
rect 4637 8128 4645 8192
rect 4325 7731 4645 8128
rect 4325 7495 4367 7731
rect 4603 7495 4645 7731
rect 4325 7104 4645 7495
rect 4325 7040 4333 7104
rect 4397 7040 4413 7104
rect 4477 7040 4493 7104
rect 4557 7040 4573 7104
rect 4637 7040 4645 7104
rect 4107 7036 4173 7037
rect 4107 6972 4108 7036
rect 4172 6972 4173 7036
rect 4107 6971 4173 6972
rect 2731 6496 2739 6560
rect 2803 6496 2819 6560
rect 2883 6496 2899 6560
rect 2963 6496 2979 6560
rect 3043 6496 3051 6560
rect 2731 6216 3051 6496
rect 2731 5980 2773 6216
rect 3009 5980 3051 6216
rect 2731 5472 3051 5980
rect 2731 5408 2739 5472
rect 2803 5408 2819 5472
rect 2883 5408 2899 5472
rect 2963 5408 2979 5472
rect 3043 5408 3051 5472
rect 2731 4384 3051 5408
rect 2731 4320 2739 4384
rect 2803 4320 2819 4384
rect 2883 4320 2899 4384
rect 2963 4320 2979 4384
rect 3043 4320 3051 4384
rect 2731 4041 3051 4320
rect 4110 4045 4170 6971
rect 4325 6016 4645 7040
rect 4325 5952 4333 6016
rect 4397 5952 4413 6016
rect 4477 5952 4493 6016
rect 4557 5952 4573 6016
rect 4637 5952 4645 6016
rect 4325 5556 4645 5952
rect 4325 5320 4367 5556
rect 4603 5320 4645 5556
rect 4325 4928 4645 5320
rect 4325 4864 4333 4928
rect 4397 4864 4413 4928
rect 4477 4864 4493 4928
rect 4557 4864 4573 4928
rect 4637 4864 4645 4928
rect 2731 3805 2773 4041
rect 3009 3805 3051 4041
rect 4107 4044 4173 4045
rect 4107 3980 4108 4044
rect 4172 3980 4173 4044
rect 4107 3979 4173 3980
rect 2731 3296 3051 3805
rect 2731 3232 2739 3296
rect 2803 3232 2819 3296
rect 2883 3232 2899 3296
rect 2963 3232 2979 3296
rect 3043 3232 3051 3296
rect 2731 2208 3051 3232
rect 2731 2144 2739 2208
rect 2803 2144 2819 2208
rect 2883 2144 2899 2208
rect 2963 2144 2979 2208
rect 3043 2144 3051 2208
rect 2731 2128 3051 2144
rect 4325 3840 4645 4864
rect 4325 3776 4333 3840
rect 4397 3776 4413 3840
rect 4477 3776 4493 3840
rect 4557 3776 4573 3840
rect 4637 3776 4645 3840
rect 4325 3381 4645 3776
rect 4325 3145 4367 3381
rect 4603 3145 4645 3381
rect 4325 2752 4645 3145
rect 4325 2688 4333 2752
rect 4397 2688 4413 2752
rect 4477 2688 4493 2752
rect 4557 2688 4573 2752
rect 4637 2688 4645 2752
rect 4325 2128 4645 2688
rect 4985 10912 5305 10928
rect 4985 10848 4993 10912
rect 5057 10848 5073 10912
rect 5137 10848 5153 10912
rect 5217 10848 5233 10912
rect 5297 10848 5305 10912
rect 4985 10566 5305 10848
rect 4985 10330 5027 10566
rect 5263 10330 5305 10566
rect 4985 9824 5305 10330
rect 4985 9760 4993 9824
rect 5057 9760 5073 9824
rect 5137 9760 5153 9824
rect 5217 9760 5233 9824
rect 5297 9760 5305 9824
rect 4985 8736 5305 9760
rect 4985 8672 4993 8736
rect 5057 8672 5073 8736
rect 5137 8672 5153 8736
rect 5217 8672 5233 8736
rect 5297 8672 5305 8736
rect 4985 8391 5305 8672
rect 4985 8155 5027 8391
rect 5263 8155 5305 8391
rect 4985 7648 5305 8155
rect 4985 7584 4993 7648
rect 5057 7584 5073 7648
rect 5137 7584 5153 7648
rect 5217 7584 5233 7648
rect 5297 7584 5305 7648
rect 4985 6560 5305 7584
rect 4985 6496 4993 6560
rect 5057 6496 5073 6560
rect 5137 6496 5153 6560
rect 5217 6496 5233 6560
rect 5297 6496 5305 6560
rect 4985 6216 5305 6496
rect 4985 5980 5027 6216
rect 5263 5980 5305 6216
rect 4985 5472 5305 5980
rect 4985 5408 4993 5472
rect 5057 5408 5073 5472
rect 5137 5408 5153 5472
rect 5217 5408 5233 5472
rect 5297 5408 5305 5472
rect 4985 4384 5305 5408
rect 4985 4320 4993 4384
rect 5057 4320 5073 4384
rect 5137 4320 5153 4384
rect 5217 4320 5233 4384
rect 5297 4320 5305 4384
rect 4985 4041 5305 4320
rect 4985 3805 5027 4041
rect 5263 3805 5305 4041
rect 4985 3296 5305 3805
rect 4985 3232 4993 3296
rect 5057 3232 5073 3296
rect 5137 3232 5153 3296
rect 5217 3232 5233 3296
rect 5297 3232 5305 3296
rect 4985 2208 5305 3232
rect 4985 2144 4993 2208
rect 5057 2144 5073 2208
rect 5137 2144 5153 2208
rect 5217 2144 5233 2208
rect 5297 2144 5305 2208
rect 4985 2128 5305 2144
rect 6579 10368 6899 10928
rect 6579 10304 6587 10368
rect 6651 10304 6667 10368
rect 6731 10304 6747 10368
rect 6811 10304 6827 10368
rect 6891 10304 6899 10368
rect 6579 9906 6899 10304
rect 6579 9670 6621 9906
rect 6857 9670 6899 9906
rect 6579 9280 6899 9670
rect 6579 9216 6587 9280
rect 6651 9216 6667 9280
rect 6731 9216 6747 9280
rect 6811 9216 6827 9280
rect 6891 9216 6899 9280
rect 6579 8192 6899 9216
rect 6579 8128 6587 8192
rect 6651 8128 6667 8192
rect 6731 8128 6747 8192
rect 6811 8128 6827 8192
rect 6891 8128 6899 8192
rect 6579 7731 6899 8128
rect 6579 7495 6621 7731
rect 6857 7495 6899 7731
rect 6579 7104 6899 7495
rect 6579 7040 6587 7104
rect 6651 7040 6667 7104
rect 6731 7040 6747 7104
rect 6811 7040 6827 7104
rect 6891 7040 6899 7104
rect 6579 6016 6899 7040
rect 6579 5952 6587 6016
rect 6651 5952 6667 6016
rect 6731 5952 6747 6016
rect 6811 5952 6827 6016
rect 6891 5952 6899 6016
rect 6579 5556 6899 5952
rect 6579 5320 6621 5556
rect 6857 5320 6899 5556
rect 6579 4928 6899 5320
rect 6579 4864 6587 4928
rect 6651 4864 6667 4928
rect 6731 4864 6747 4928
rect 6811 4864 6827 4928
rect 6891 4864 6899 4928
rect 6579 3840 6899 4864
rect 6579 3776 6587 3840
rect 6651 3776 6667 3840
rect 6731 3776 6747 3840
rect 6811 3776 6827 3840
rect 6891 3776 6899 3840
rect 6579 3381 6899 3776
rect 6579 3145 6621 3381
rect 6857 3145 6899 3381
rect 6579 2752 6899 3145
rect 6579 2688 6587 2752
rect 6651 2688 6667 2752
rect 6731 2688 6747 2752
rect 6811 2688 6827 2752
rect 6891 2688 6899 2752
rect 6579 2128 6899 2688
rect 7239 10912 7559 10928
rect 7239 10848 7247 10912
rect 7311 10848 7327 10912
rect 7391 10848 7407 10912
rect 7471 10848 7487 10912
rect 7551 10848 7559 10912
rect 7239 10566 7559 10848
rect 7239 10330 7281 10566
rect 7517 10330 7559 10566
rect 7239 9824 7559 10330
rect 7239 9760 7247 9824
rect 7311 9760 7327 9824
rect 7391 9760 7407 9824
rect 7471 9760 7487 9824
rect 7551 9760 7559 9824
rect 7239 8736 7559 9760
rect 7239 8672 7247 8736
rect 7311 8672 7327 8736
rect 7391 8672 7407 8736
rect 7471 8672 7487 8736
rect 7551 8672 7559 8736
rect 7239 8391 7559 8672
rect 7239 8155 7281 8391
rect 7517 8155 7559 8391
rect 7239 7648 7559 8155
rect 7239 7584 7247 7648
rect 7311 7584 7327 7648
rect 7391 7584 7407 7648
rect 7471 7584 7487 7648
rect 7551 7584 7559 7648
rect 7239 6560 7559 7584
rect 7239 6496 7247 6560
rect 7311 6496 7327 6560
rect 7391 6496 7407 6560
rect 7471 6496 7487 6560
rect 7551 6496 7559 6560
rect 7239 6216 7559 6496
rect 7239 5980 7281 6216
rect 7517 5980 7559 6216
rect 7239 5472 7559 5980
rect 7239 5408 7247 5472
rect 7311 5408 7327 5472
rect 7391 5408 7407 5472
rect 7471 5408 7487 5472
rect 7551 5408 7559 5472
rect 7239 4384 7559 5408
rect 7239 4320 7247 4384
rect 7311 4320 7327 4384
rect 7391 4320 7407 4384
rect 7471 4320 7487 4384
rect 7551 4320 7559 4384
rect 7239 4041 7559 4320
rect 7239 3805 7281 4041
rect 7517 3805 7559 4041
rect 7239 3296 7559 3805
rect 7239 3232 7247 3296
rect 7311 3232 7327 3296
rect 7391 3232 7407 3296
rect 7471 3232 7487 3296
rect 7551 3232 7559 3296
rect 7239 2208 7559 3232
rect 7239 2144 7247 2208
rect 7311 2144 7327 2208
rect 7391 2144 7407 2208
rect 7471 2144 7487 2208
rect 7551 2144 7559 2208
rect 7239 2128 7559 2144
rect 8833 10368 9153 10928
rect 8833 10304 8841 10368
rect 8905 10304 8921 10368
rect 8985 10304 9001 10368
rect 9065 10304 9081 10368
rect 9145 10304 9153 10368
rect 8833 9906 9153 10304
rect 8833 9670 8875 9906
rect 9111 9670 9153 9906
rect 8833 9280 9153 9670
rect 8833 9216 8841 9280
rect 8905 9216 8921 9280
rect 8985 9216 9001 9280
rect 9065 9216 9081 9280
rect 9145 9216 9153 9280
rect 8833 8192 9153 9216
rect 8833 8128 8841 8192
rect 8905 8128 8921 8192
rect 8985 8128 9001 8192
rect 9065 8128 9081 8192
rect 9145 8128 9153 8192
rect 8833 7731 9153 8128
rect 8833 7495 8875 7731
rect 9111 7495 9153 7731
rect 8833 7104 9153 7495
rect 8833 7040 8841 7104
rect 8905 7040 8921 7104
rect 8985 7040 9001 7104
rect 9065 7040 9081 7104
rect 9145 7040 9153 7104
rect 8833 6016 9153 7040
rect 8833 5952 8841 6016
rect 8905 5952 8921 6016
rect 8985 5952 9001 6016
rect 9065 5952 9081 6016
rect 9145 5952 9153 6016
rect 8833 5556 9153 5952
rect 8833 5320 8875 5556
rect 9111 5320 9153 5556
rect 8833 4928 9153 5320
rect 8833 4864 8841 4928
rect 8905 4864 8921 4928
rect 8985 4864 9001 4928
rect 9065 4864 9081 4928
rect 9145 4864 9153 4928
rect 8833 3840 9153 4864
rect 8833 3776 8841 3840
rect 8905 3776 8921 3840
rect 8985 3776 9001 3840
rect 9065 3776 9081 3840
rect 9145 3776 9153 3840
rect 8833 3381 9153 3776
rect 8833 3145 8875 3381
rect 9111 3145 9153 3381
rect 8833 2752 9153 3145
rect 8833 2688 8841 2752
rect 8905 2688 8921 2752
rect 8985 2688 9001 2752
rect 9065 2688 9081 2752
rect 9145 2688 9153 2752
rect 8833 2128 9153 2688
rect 9493 10912 9813 10928
rect 9493 10848 9501 10912
rect 9565 10848 9581 10912
rect 9645 10848 9661 10912
rect 9725 10848 9741 10912
rect 9805 10848 9813 10912
rect 9493 10566 9813 10848
rect 9493 10330 9535 10566
rect 9771 10330 9813 10566
rect 9493 9824 9813 10330
rect 9493 9760 9501 9824
rect 9565 9760 9581 9824
rect 9645 9760 9661 9824
rect 9725 9760 9741 9824
rect 9805 9760 9813 9824
rect 9493 8736 9813 9760
rect 9493 8672 9501 8736
rect 9565 8672 9581 8736
rect 9645 8672 9661 8736
rect 9725 8672 9741 8736
rect 9805 8672 9813 8736
rect 9493 8391 9813 8672
rect 9493 8155 9535 8391
rect 9771 8155 9813 8391
rect 9493 7648 9813 8155
rect 9493 7584 9501 7648
rect 9565 7584 9581 7648
rect 9645 7584 9661 7648
rect 9725 7584 9741 7648
rect 9805 7584 9813 7648
rect 9493 6560 9813 7584
rect 9493 6496 9501 6560
rect 9565 6496 9581 6560
rect 9645 6496 9661 6560
rect 9725 6496 9741 6560
rect 9805 6496 9813 6560
rect 9493 6216 9813 6496
rect 9493 5980 9535 6216
rect 9771 5980 9813 6216
rect 9493 5472 9813 5980
rect 9493 5408 9501 5472
rect 9565 5408 9581 5472
rect 9645 5408 9661 5472
rect 9725 5408 9741 5472
rect 9805 5408 9813 5472
rect 9493 4384 9813 5408
rect 9493 4320 9501 4384
rect 9565 4320 9581 4384
rect 9645 4320 9661 4384
rect 9725 4320 9741 4384
rect 9805 4320 9813 4384
rect 9493 4041 9813 4320
rect 9493 3805 9535 4041
rect 9771 3805 9813 4041
rect 9493 3296 9813 3805
rect 9493 3232 9501 3296
rect 9565 3232 9581 3296
rect 9645 3232 9661 3296
rect 9725 3232 9741 3296
rect 9805 3232 9813 3296
rect 9493 2208 9813 3232
rect 9493 2144 9501 2208
rect 9565 2144 9581 2208
rect 9645 2144 9661 2208
rect 9725 2144 9741 2208
rect 9805 2144 9813 2208
rect 9493 2128 9813 2144
<< via4 >>
rect 2113 9670 2349 9906
rect 2113 7495 2349 7731
rect 2113 5320 2349 5556
rect 2113 3145 2349 3381
rect 2773 10330 3009 10566
rect 2773 8155 3009 8391
rect 4367 9670 4603 9906
rect 4367 7495 4603 7731
rect 2773 5980 3009 6216
rect 4367 5320 4603 5556
rect 2773 3805 3009 4041
rect 4367 3145 4603 3381
rect 5027 10330 5263 10566
rect 5027 8155 5263 8391
rect 5027 5980 5263 6216
rect 5027 3805 5263 4041
rect 6621 9670 6857 9906
rect 6621 7495 6857 7731
rect 6621 5320 6857 5556
rect 6621 3145 6857 3381
rect 7281 10330 7517 10566
rect 7281 8155 7517 8391
rect 7281 5980 7517 6216
rect 7281 3805 7517 4041
rect 8875 9670 9111 9906
rect 8875 7495 9111 7731
rect 8875 5320 9111 5556
rect 8875 3145 9111 3381
rect 9535 10330 9771 10566
rect 9535 8155 9771 8391
rect 9535 5980 9771 6216
rect 9535 3805 9771 4041
<< metal5 >>
rect 1056 10566 10168 10608
rect 1056 10330 2773 10566
rect 3009 10330 5027 10566
rect 5263 10330 7281 10566
rect 7517 10330 9535 10566
rect 9771 10330 10168 10566
rect 1056 10288 10168 10330
rect 1056 9906 10168 9948
rect 1056 9670 2113 9906
rect 2349 9670 4367 9906
rect 4603 9670 6621 9906
rect 6857 9670 8875 9906
rect 9111 9670 10168 9906
rect 1056 9628 10168 9670
rect 1056 8391 10168 8433
rect 1056 8155 2773 8391
rect 3009 8155 5027 8391
rect 5263 8155 7281 8391
rect 7517 8155 9535 8391
rect 9771 8155 10168 8391
rect 1056 8113 10168 8155
rect 1056 7731 10168 7773
rect 1056 7495 2113 7731
rect 2349 7495 4367 7731
rect 4603 7495 6621 7731
rect 6857 7495 8875 7731
rect 9111 7495 10168 7731
rect 1056 7453 10168 7495
rect 1056 6216 10168 6258
rect 1056 5980 2773 6216
rect 3009 5980 5027 6216
rect 5263 5980 7281 6216
rect 7517 5980 9535 6216
rect 9771 5980 10168 6216
rect 1056 5938 10168 5980
rect 1056 5556 10168 5598
rect 1056 5320 2113 5556
rect 2349 5320 4367 5556
rect 4603 5320 6621 5556
rect 6857 5320 8875 5556
rect 9111 5320 10168 5556
rect 1056 5278 10168 5320
rect 1056 4041 10168 4083
rect 1056 3805 2773 4041
rect 3009 3805 5027 4041
rect 5263 3805 7281 4041
rect 7517 3805 9535 4041
rect 9771 3805 10168 4041
rect 1056 3763 10168 3805
rect 1056 3381 10168 3423
rect 1056 3145 2113 3381
rect 2349 3145 4367 3381
rect 4603 3145 6621 3381
rect 6857 3145 8875 3381
rect 9111 3145 10168 3381
rect 1056 3103 10168 3145
use sky130_fd_sc_hd__or2_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5520 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _22_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4416 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _23_
timestamp 1723858470
transform 1 0 4140 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _24_
timestamp 1723858470
transform 1 0 4692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _25_
timestamp 1723858470
transform 1 0 4600 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _26_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 4876 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _27_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5152 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _28_
timestamp 1723858470
transform -1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _29_
timestamp 1723858470
transform -1 0 5888 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _30_
timestamp 1723858470
transform -1 0 4876 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _31_
timestamp 1723858470
transform -1 0 8648 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _32_
timestamp 1723858470
transform -1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _33_
timestamp 1723858470
transform -1 0 8280 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _34_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 8648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _35_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _36_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _37_
timestamp 1723858470
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6992 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6440 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _40_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 6348 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5152 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _42_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5060 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _43_
timestamp 1723858470
transform -1 0 5428 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _44_
timestamp 1723858470
transform -1 0 4784 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _45_
timestamp 1723858470
transform 1 0 7636 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _46_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 5612 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _47_
timestamp 1723858470
transform -1 0 3220 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _48_
timestamp 1723858470
transform -1 0 3220 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _49_
timestamp 1723858470
transform 1 0 6992 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _50_
timestamp 1723858470
transform 1 0 6992 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _51_
timestamp 1723858470
transform -1 0 3220 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _52_
timestamp 1723858470
transform -1 0 8464 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _53_
timestamp 1723858470
transform -1 0 5520 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _54_
timestamp 1723858470
transform 1 0 1840 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _55_
timestamp 1723858470
transform 1 0 6532 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _56_
timestamp 1723858470
transform 1 0 3404 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _57_
timestamp 1723858470
transform -1 0 3680 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _58_
timestamp 1723858470
transform -1 0 6900 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _59_
timestamp 1723858470
transform 1 0 6808 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _60_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6900 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5152 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1723858470
transform -1 0 3772 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1723858470
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout17 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 4324 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5244 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_41
timestamp 1723858470
transform 1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1723858470
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1723858470
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_85
timestamp 1723858470
transform 1 0 8924 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_91
timestamp 1723858470
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_49
timestamp 1723858470
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1723858470
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_61
timestamp 1723858470
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_82
timestamp 1723858470
transform 1 0 8648 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_90
timestamp 1723858470
transform 1 0 9384 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1723858470
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1723858470
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1723858470
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1723858470
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1723858470
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_53
timestamp 1723858470
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_61
timestamp 1723858470
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1723858470
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_93
timestamp 1723858470
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1723858470
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1723858470
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1723858470
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1723858470
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1723858470
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1723858470
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1723858470
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1723858470
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1723858470
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_93
timestamp 1723858470
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1723858470
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1723858470
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1723858470
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1723858470
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1723858470
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1723858470
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_68
timestamp 1723858470
transform 1 0 7360 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_72
timestamp 1723858470
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1723858470
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_93
timestamp 1723858470
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_3
timestamp 1723858470
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_7
timestamp 1723858470
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_48
timestamp 1723858470
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1723858470
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_82
timestamp 1723858470
transform 1 0 8648 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_94
timestamp 1723858470
transform 1 0 9752 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 1723858470
transform 1 0 1656 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1723858470
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1723858470
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_35
timestamp 1723858470
transform 1 0 4324 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_50
timestamp 1723858470
transform 1 0 5704 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_62
timestamp 1723858470
transform 1 0 6808 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_88
timestamp 1723858470
transform 1 0 9200 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1723858470
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1723858470
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_27
timestamp 1723858470
transform 1 0 3588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_49
timestamp 1723858470
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1723858470
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1723858470
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_72
timestamp 1723858470
transform 1 0 7728 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_82
timestamp 1723858470
transform 1 0 8648 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_94
timestamp 1723858470
transform 1 0 9752 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1723858470
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1723858470
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1723858470
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1723858470
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_37
timestamp 1723858470
transform 1 0 4508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_64
timestamp 1723858470
transform 1 0 6992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_76
timestamp 1723858470
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1723858470
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_93
timestamp 1723858470
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1723858470
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 1723858470
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_49
timestamp 1723858470
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1723858470
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1723858470
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_69
timestamp 1723858470
transform 1 0 7452 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_77
timestamp 1723858470
transform 1 0 8188 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_87
timestamp 1723858470
transform 1 0 9108 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1723858470
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1723858470
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1723858470
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1723858470
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_57
timestamp 1723858470
transform 1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_79
timestamp 1723858470
transform 1 0 8372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1723858470
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1723858470
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_93
timestamp 1723858470
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_23
timestamp 1723858470
transform 1 0 3220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49
timestamp 1723858470
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1723858470
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_57
timestamp 1723858470
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_80
timestamp 1723858470
transform 1 0 8464 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_92
timestamp 1723858470
transform 1 0 9568 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1723858470
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1723858470
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1723858470
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1723858470
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1723858470
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_53
timestamp 1723858470
transform 1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_57
timestamp 1723858470
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_66
timestamp 1723858470
transform 1 0 7176 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_78
timestamp 1723858470
transform 1 0 8280 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_85
timestamp 1723858470
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_91
timestamp 1723858470
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_23
timestamp 1723858470
transform 1 0 3220 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_52
timestamp 1723858470
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1723858470
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1723858470
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1723858470
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_93
timestamp 1723858470
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1723858470
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_7
timestamp 1723858470
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1723858470
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1723858470
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_93
timestamp 1723858470
transform 1 0 9660 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_12
timestamp 1723858470
transform 1 0 2208 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_24
timestamp 1723858470
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_29
timestamp 1723858470
transform 1 0 3772 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_34
timestamp 1723858470
transform 1 0 4232 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_42
timestamp 1723858470
transform 1 0 4968 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_48
timestamp 1723858470
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1723858470
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 1723858470
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1723858470
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_81
timestamp 1723858470
transform 1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_85
timestamp 1723858470
transform 1 0 8924 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform -1 0 7176 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1723858470
transform -1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1723858470
transform 1 0 8372 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9568 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1723858470
transform 1 0 9568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1723858470
transform -1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1723858470
transform 1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1723858470
transform 1 0 3956 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1723858470
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1723858470
transform 1 0 9292 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1723858470
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1723858470
transform 1 0 9568 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 9476 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 1723858470
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1723858470
transform 1 0 5060 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1723858470
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1723858470
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 1723858470
transform 1 0 9292 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1723858470
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1723858470
transform -1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1723858470
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1723858470
transform -1 0 10120 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1723858470
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1723858470
transform -1 0 10120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1723858470
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1723858470
transform -1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1723858470
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1723858470
transform -1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1723858470
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1723858470
transform -1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1723858470
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1723858470
transform -1 0 10120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1723858470
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1723858470
transform -1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1723858470
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1723858470
transform -1 0 10120 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1723858470
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1723858470
transform -1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1723858470
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1723858470
transform -1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1723858470
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1723858470
transform -1 0 10120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1723858470
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1723858470
transform -1 0 10120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1723858470
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1723858470
transform -1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1723858470
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1723858470
transform -1 0 10120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1723858470
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1723858470
transform -1 0 10120 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1723858470
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1723858470
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1723858470
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1723858470
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1723858470
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1723858470
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1723858470
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1723858470
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1723858470
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1723858470
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1723858470
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1723858470
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1723858470
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1723858470
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1723858470
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1723858470
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1723858470
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1723858470
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1723858470
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1723858470
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1723858470
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1723858470
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1723858470
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1723858470
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1723858470
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1723858470
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1723858470
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
<< labels >>
flabel metal4 s 2731 2128 3051 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4985 2128 5305 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7239 2128 7559 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 9493 2128 9813 10928 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3763 10168 4083 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5938 10168 6258 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8113 10168 8433 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 10288 10168 10608 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2071 2128 2391 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 4325 2128 4645 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6579 2128 6899 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8833 2128 9153 10928 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3103 10168 3423 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5278 10168 5598 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7453 10168 7773 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 9628 10168 9948 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 10495 8848 11295 8968 0 FreeSans 480 0 0 0 a_in[0]
port 2 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 a_in[1]
port 3 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 a_in[2]
port 4 nsew signal input
flabel metal2 s 7102 12639 7158 13439 0 FreeSans 224 90 0 0 a_in[3]
port 5 nsew signal input
flabel metal2 s 3882 12639 3938 13439 0 FreeSans 224 90 0 0 b_in[0]
port 6 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 b_in[1]
port 7 nsew signal input
flabel metal3 s 10495 11568 11295 11688 0 FreeSans 480 0 0 0 b_in[2]
port 8 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 b_in[3]
port 9 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 clk
port 10 nsew signal input
flabel metal3 s 10495 2728 11295 2848 0 FreeSans 480 0 0 0 cout_out
port 11 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 ovf_out
port 12 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 rst_n
port 13 nsew signal input
flabel metal2 s 9678 12639 9734 13439 0 FreeSans 224 90 0 0 sub_in
port 14 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 y_out[0]
port 15 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 y_out[1]
port 16 nsew signal tristate
flabel metal2 s 1306 12639 1362 13439 0 FreeSans 224 90 0 0 y_out[2]
port 17 nsew signal tristate
flabel metal3 s 10495 5448 11295 5568 0 FreeSans 480 0 0 0 y_out[3]
port 18 nsew signal tristate
rlabel metal1 5612 10880 5612 10880 0 VGND
rlabel metal1 5612 10336 5612 10336 0 VPWR
rlabel metal1 5336 10438 5336 10438 0 _00_
rlabel metal1 5336 9894 5336 9894 0 _01_
rlabel metal1 4370 9690 4370 9690 0 _02_
rlabel metal1 4784 6358 4784 6358 0 _03_
rlabel metal1 5106 6222 5106 6222 0 _04_
rlabel metal1 5014 6766 5014 6766 0 _05_
rlabel metal1 4922 7412 4922 7412 0 _06_
rlabel metal1 5290 6970 5290 6970 0 _07_
rlabel metal1 4370 9520 4370 9520 0 _08_
rlabel metal1 5382 9350 5382 9350 0 _09_
rlabel metal1 7038 5134 7038 5134 0 _10_
rlabel via1 8234 6086 8234 6086 0 _11_
rlabel metal1 8326 6222 8326 6222 0 _12_
rlabel metal1 7498 6256 7498 6256 0 _13_
rlabel metal1 7774 6290 7774 6290 0 _14_
rlabel metal1 7590 5134 7590 5134 0 _15_
rlabel metal1 7728 4794 7728 4794 0 _16_
rlabel metal2 7222 4998 7222 4998 0 _17_
rlabel metal1 4738 6834 4738 6834 0 _18_
rlabel metal1 4738 9690 4738 9690 0 _19_
rlabel metal1 9982 8942 9982 8942 0 a_in[0]
rlabel metal2 10994 1588 10994 1588 0 a_in[1]
rlabel metal3 1326 11628 1326 11628 0 a_in[2]
rlabel metal1 7268 10642 7268 10642 0 a_in[3]
rlabel metal1 6670 8296 6670 8296 0 a_r\[0\]
rlabel metal2 4830 5712 4830 5712 0 a_r\[1\]
rlabel metal1 4646 10676 4646 10676 0 a_r\[2\]
rlabel metal1 8372 7378 8372 7378 0 a_r\[3\]
rlabel metal1 4048 10642 4048 10642 0 b_in[0]
rlabel metal2 46 1520 46 1520 0 b_in[1]
rlabel metal1 9430 10642 9430 10642 0 b_in[2]
rlabel metal2 8418 1588 8418 1588 0 b_in[3]
rlabel metal1 5336 7922 5336 7922 0 b_r\[0\]
rlabel metal1 4738 5644 4738 5644 0 b_r\[1\]
rlabel metal1 5198 10234 5198 10234 0 b_r\[2\]
rlabel metal2 8602 4182 8602 4182 0 b_r\[3\]
rlabel metal2 2622 2115 2622 2115 0 clk
rlabel metal1 4278 7378 4278 7378 0 clknet_0_clk
rlabel metal1 3036 2482 3036 2482 0 clknet_1_0__leaf_clk
rlabel metal1 6578 7990 6578 7990 0 clknet_1_1__leaf_clk
rlabel via2 9706 2805 9706 2805 0 cout_out
rlabel metal1 8510 8534 8510 8534 0 net1
rlabel metal1 8418 10098 8418 10098 0 net10
rlabel metal1 9154 3026 9154 3026 0 net11
rlabel metal1 1472 2618 1472 2618 0 net12
rlabel metal1 4968 2414 4968 2414 0 net13
rlabel metal1 1472 8602 1472 8602 0 net14
rlabel metal1 1472 9690 1472 9690 0 net15
rlabel metal1 9108 5610 9108 5610 0 net16
rlabel metal2 2438 3570 2438 3570 0 net17
rlabel metal1 4370 9962 4370 9962 0 net18
rlabel metal1 6210 7854 6210 7854 0 net19
rlabel metal1 9154 2618 9154 2618 0 net2
rlabel metal1 5336 3094 5336 3094 0 net20
rlabel metal1 8694 6358 8694 6358 0 net21
rlabel metal1 2060 10234 2060 10234 0 net3
rlabel metal1 6624 7786 6624 7786 0 net4
rlabel metal1 3864 8534 3864 8534 0 net5
rlabel metal1 3312 2618 3312 2618 0 net6
rlabel metal1 7967 10234 7967 10234 0 net7
rlabel metal1 7820 2958 7820 2958 0 net8
rlabel metal1 1610 5576 1610 5576 0 net9
rlabel metal1 3128 2346 3128 2346 0 ovf
rlabel metal3 820 2788 820 2788 0 ovf_out
rlabel metal3 1050 5508 1050 5508 0 rst_n
rlabel metal1 9844 10642 9844 10642 0 sub_in
rlabel metal1 5382 7786 5382 7786 0 sub_r
rlabel metal1 5704 5746 5704 5746 0 sum\[0\]
rlabel metal1 4324 7514 4324 7514 0 sum\[1\]
rlabel metal1 3542 9622 3542 9622 0 sum\[2\]
rlabel metal2 7038 5440 7038 5440 0 sum\[3\]
rlabel metal1 7498 3570 7498 3570 0 sum\[4\]
rlabel metal2 5198 959 5198 959 0 y_out[0]
rlabel metal3 820 8908 820 8908 0 y_out[1]
rlabel metal1 1472 10778 1472 10778 0 y_out[2]
rlabel metal1 9890 5542 9890 5542 0 y_out[3]
<< properties >>
string FIXED_BBOX 0 0 11295 13439
<< end >>
