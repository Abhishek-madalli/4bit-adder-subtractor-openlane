VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO addsub4_top
  CLASS BLOCK ;
  FOREIGN addsub4_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 56.475 BY 67.195 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.655 10.640 15.255 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.925 10.640 26.525 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.195 10.640 37.795 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.465 10.640 49.065 54.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.815 50.840 20.415 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 29.690 50.840 31.290 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 40.565 50.840 42.165 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 51.440 50.840 53.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.355 10.640 11.955 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.625 10.640 23.225 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.895 10.640 34.495 54.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.165 10.640 45.765 54.640 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 15.515 50.840 17.115 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.390 50.840 27.990 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 37.265 50.840 38.865 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 48.140 50.840 49.740 ;
    END
  END VPWR
  PIN a_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 52.475 44.240 56.475 44.840 ;
    END
  END a_in[0]
  PIN a_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END a_in[1]
  PIN a_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END a_in[2]
  PIN a_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 63.195 35.790 67.195 ;
    END
  END a_in[3]
  PIN b_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 63.195 19.690 67.195 ;
    END
  END b_in[0]
  PIN b_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END b_in[1]
  PIN b_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 52.475 57.840 56.475 58.440 ;
    END
  END b_in[2]
  PIN b_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END b_in[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END clk
  PIN cout_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 52.475 13.640 56.475 14.240 ;
    END
  END cout_out
  PIN ovf_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END ovf_out
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END rst_n
  PIN sub_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 63.195 48.670 67.195 ;
    END
  END sub_in
  PIN y_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END y_out[0]
  PIN y_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END y_out[1]
  PIN y_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 6.530 63.195 6.810 67.195 ;
    END
  END y_out[2]
  PIN y_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 52.475 27.240 56.475 27.840 ;
    END
  END y_out[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 50.600 54.485 ;
      LAYER met1 ;
        RECT 0.070 10.640 55.130 54.640 ;
      LAYER met2 ;
        RECT 0.100 62.915 6.250 63.195 ;
        RECT 7.090 62.915 19.130 63.195 ;
        RECT 19.970 62.915 35.230 63.195 ;
        RECT 36.070 62.915 48.110 63.195 ;
        RECT 48.950 62.915 55.100 63.195 ;
        RECT 0.100 4.280 55.100 62.915 ;
        RECT 0.650 4.000 12.690 4.280 ;
        RECT 13.530 4.000 25.570 4.280 ;
        RECT 26.410 4.000 41.670 4.280 ;
        RECT 42.510 4.000 54.550 4.280 ;
      LAYER met3 ;
        RECT 4.400 57.440 52.075 58.305 ;
        RECT 4.000 45.240 52.475 57.440 ;
        RECT 4.400 43.840 52.075 45.240 ;
        RECT 4.000 28.240 52.475 43.840 ;
        RECT 4.400 26.840 52.075 28.240 ;
        RECT 4.000 14.640 52.475 26.840 ;
        RECT 4.400 13.240 52.075 14.640 ;
        RECT 4.000 10.715 52.475 13.240 ;
      LAYER met4 ;
        RECT 20.535 19.895 20.865 35.185 ;
  END
END addsub4_top
END LIBRARY

