magic
tech sky130A
magscale 1 2
timestamp 1755103507
<< obsli1 >>
rect 1104 2159 10120 10897
<< obsm1 >>
rect 14 2128 11026 10928
<< metal2 >>
rect 1306 12639 1362 13439
rect 3882 12639 3938 13439
rect 7102 12639 7158 13439
rect 9678 12639 9734 13439
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 8390 0 8446 800
rect 10966 0 11022 800
<< obsm2 >>
rect 20 12583 1250 12639
rect 1418 12583 3826 12639
rect 3994 12583 7046 12639
rect 7214 12583 9622 12639
rect 9790 12583 11020 12639
rect 20 856 11020 12583
rect 130 800 2538 856
rect 2706 800 5114 856
rect 5282 800 8334 856
rect 8502 800 10910 856
<< metal3 >>
rect 0 11568 800 11688
rect 10495 11568 11295 11688
rect 0 8848 800 8968
rect 10495 8848 11295 8968
rect 0 5448 800 5568
rect 10495 5448 11295 5568
rect 0 2728 800 2848
rect 10495 2728 11295 2848
<< obsm3 >>
rect 880 11488 10415 11661
rect 800 9048 10495 11488
rect 880 8768 10415 9048
rect 800 5648 10495 8768
rect 880 5368 10415 5648
rect 800 2928 10495 5368
rect 880 2648 10415 2928
rect 800 2143 10495 2648
<< metal4 >>
rect 2071 2128 2391 10928
rect 2731 2128 3051 10928
rect 4325 2128 4645 10928
rect 4985 2128 5305 10928
rect 6579 2128 6899 10928
rect 7239 2128 7559 10928
rect 8833 2128 9153 10928
rect 9493 2128 9813 10928
<< obsm4 >>
rect 4107 3979 4173 7037
<< metal5 >>
rect 1056 10288 10168 10608
rect 1056 9628 10168 9948
rect 1056 8113 10168 8433
rect 1056 7453 10168 7773
rect 1056 5938 10168 6258
rect 1056 5278 10168 5598
rect 1056 3763 10168 4083
rect 1056 3103 10168 3423
<< labels >>
rlabel metal4 s 2731 2128 3051 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4985 2128 5305 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7239 2128 7559 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 9493 2128 9813 10928 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3763 10168 4083 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5938 10168 6258 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8113 10168 8433 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 10288 10168 10608 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2071 2128 2391 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4325 2128 4645 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 6579 2128 6899 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 8833 2128 9153 10928 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3103 10168 3423 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5278 10168 5598 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7453 10168 7773 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 9628 10168 9948 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 10495 8848 11295 8968 6 a_in[0]
port 3 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 a_in[1]
port 4 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 a_in[2]
port 5 nsew signal input
rlabel metal2 s 7102 12639 7158 13439 6 a_in[3]
port 6 nsew signal input
rlabel metal2 s 3882 12639 3938 13439 6 b_in[0]
port 7 nsew signal input
rlabel metal2 s 18 0 74 800 6 b_in[1]
port 8 nsew signal input
rlabel metal3 s 10495 11568 11295 11688 6 b_in[2]
port 9 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 b_in[3]
port 10 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 clk
port 11 nsew signal input
rlabel metal3 s 10495 2728 11295 2848 6 cout_out
port 12 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 ovf_out
port 13 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 rst_n
port 14 nsew signal input
rlabel metal2 s 9678 12639 9734 13439 6 sub_in
port 15 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 y_out[0]
port 16 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 y_out[1]
port 17 nsew signal output
rlabel metal2 s 1306 12639 1362 13439 6 y_out[2]
port 18 nsew signal output
rlabel metal3 s 10495 5448 11295 5568 6 y_out[3]
port 19 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 11295 13439
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 370392
string GDS_FILE /openlane/designs/addsub4/runs/run1/results/signoff/addsub4_top.magic.gds
string GDS_START 160480
<< end >>

